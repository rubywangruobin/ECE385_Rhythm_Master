module who_win(input Reset, frame_clk, 
						input logic [7:0] keycode,
						 input [13:0] total_Score, total_Score_1,
						 output logic [2249:0] tie_graph,
						 output logic [2374:0] win_graph,
						 output logic [1:0] winner);
	logic [11:0] counter;
	 enum logic [3:0] {Halted, Normal, End} State, Next_state;
	 logic finish_on;
	 always_ff @ (posedge frame_clk )
    begin
		if(Reset)
		begin
			State <= Halted;
		end	
		else if(State == Halted)
		begin
			counter = 0;
			winner = 2'b00;
			State <= Next_state;
		end
		else if(State == Normal)
			begin
				if(counter <3500)
					counter = counter + 1;
				else
					begin
						if(total_Score > total_Score_1)
							winner = 2'b01;
						else if(total_Score < total_Score_1)
							winner = 2'b10;
						else
							winner= 2'b00;
					end
				State <= Next_state;
			end
		else
			State <= Next_state;
    end
	 
	 always_comb
	 begin
		Next_state = State;
		finish_on = 1'b0;
		unique case(State)
			Halted:
			begin
				finish_on = 1'b0;
				if(keycode == 8'h2c)
					Next_state = Normal;
			end
			Normal:
				begin
				if(counter < 3500)
					Next_state = Normal;
				else
					Next_state = End;
				end
			End:
				begin
				finish_on = 1;
				if(keycode == 8'h01)
					Next_state = Halted;
				end
		endcase
					
	 end
	 always_comb
	 begin
		tie_graph <= 1'b0;
		win_graph <= 1'b0;
		if(finish_on == 1)
		begin
		case(winner)
			2'b00:
				begin
					tie_graph[338] <= 1'b1;
tie_graph[339] <= 1'b1;
tie_graph[360] <= 1'b1;
tie_graph[361] <= 1'b1;
tie_graph[374] <= 1'b1;
tie_graph[375] <= 1'b1;
tie_graph[414] <= 1'b1;
tie_graph[415] <= 1'b1;
tie_graph[416] <= 1'b1;
tie_graph[417] <= 1'b1;
tie_graph[418] <= 1'b1;
tie_graph[419] <= 1'b1;
tie_graph[420] <= 1'b1;
tie_graph[421] <= 1'b1;
tie_graph[422] <= 1'b1;
tie_graph[423] <= 1'b1;
tie_graph[424] <= 1'b1;
tie_graph[425] <= 1'b1;
tie_graph[428] <= 1'b1;
tie_graph[429] <= 1'b1;
tie_graph[447] <= 1'b1;
tie_graph[448] <= 1'b1;
tie_graph[450] <= 1'b1;
tie_graph[451] <= 1'b1;
tie_graph[457] <= 1'b1;
tie_graph[458] <= 1'b1;
tie_graph[464] <= 1'b1;
tie_graph[465] <= 1'b1;
tie_graph[504] <= 1'b1;
tie_graph[505] <= 1'b1;
tie_graph[506] <= 1'b1;
tie_graph[507] <= 1'b1;
tie_graph[508] <= 1'b1;
tie_graph[509] <= 1'b1;
tie_graph[510] <= 1'b1;
tie_graph[511] <= 1'b1;
tie_graph[512] <= 1'b1;
tie_graph[513] <= 1'b1;
tie_graph[514] <= 1'b1;
tie_graph[515] <= 1'b1;
tie_graph[537] <= 1'b1;
tie_graph[538] <= 1'b1;
tie_graph[540] <= 1'b1;
tie_graph[541] <= 1'b1;
tie_graph[547] <= 1'b1;
tie_graph[548] <= 1'b1;
tie_graph[554] <= 1'b1;
tie_graph[555] <= 1'b1;
tie_graph[599] <= 1'b1;
tie_graph[600] <= 1'b1;
tie_graph[627] <= 1'b1;
tie_graph[628] <= 1'b1;
tie_graph[630] <= 1'b1;
tie_graph[631] <= 1'b1;
tie_graph[637] <= 1'b1;
tie_graph[638] <= 1'b1;
tie_graph[644] <= 1'b1;
tie_graph[645] <= 1'b1;
tie_graph[689] <= 1'b1;
tie_graph[690] <= 1'b1;
tie_graph[717] <= 1'b1;
tie_graph[718] <= 1'b1;
tie_graph[720] <= 1'b1;
tie_graph[721] <= 1'b1;
tie_graph[725] <= 1'b1;
tie_graph[726] <= 1'b1;
tie_graph[727] <= 1'b1;
tie_graph[728] <= 1'b1;
tie_graph[729] <= 1'b1;
tie_graph[730] <= 1'b1;
tie_graph[731] <= 1'b1;
tie_graph[734] <= 1'b1;
tie_graph[735] <= 1'b1;
tie_graph[743] <= 1'b1;
tie_graph[744] <= 1'b1;
tie_graph[758] <= 1'b1;
tie_graph[759] <= 1'b1;
tie_graph[760] <= 1'b1;
tie_graph[761] <= 1'b1;
tie_graph[762] <= 1'b1;
tie_graph[779] <= 1'b1;
tie_graph[780] <= 1'b1;
tie_graph[796] <= 1'b1;
tie_graph[797] <= 1'b1;
tie_graph[798] <= 1'b1;
tie_graph[799] <= 1'b1;
tie_graph[800] <= 1'b1;
tie_graph[807] <= 1'b1;
tie_graph[808] <= 1'b1;
tie_graph[810] <= 1'b1;
tie_graph[811] <= 1'b1;
tie_graph[815] <= 1'b1;
tie_graph[816] <= 1'b1;
tie_graph[817] <= 1'b1;
tie_graph[818] <= 1'b1;
tie_graph[819] <= 1'b1;
tie_graph[820] <= 1'b1;
tie_graph[821] <= 1'b1;
tie_graph[831] <= 1'b1;
tie_graph[832] <= 1'b1;
tie_graph[833] <= 1'b1;
tie_graph[834] <= 1'b1;
tie_graph[835] <= 1'b1;
tie_graph[836] <= 1'b1;
tie_graph[847] <= 1'b1;
tie_graph[848] <= 1'b1;
tie_graph[849] <= 1'b1;
tie_graph[850] <= 1'b1;
tie_graph[851] <= 1'b1;
tie_graph[852] <= 1'b1;
tie_graph[853] <= 1'b1;
tie_graph[869] <= 1'b1;
tie_graph[870] <= 1'b1;
tie_graph[878] <= 1'b1;
tie_graph[879] <= 1'b1;
tie_graph[885] <= 1'b1;
tie_graph[886] <= 1'b1;
tie_graph[887] <= 1'b1;
tie_graph[889] <= 1'b1;
tie_graph[890] <= 1'b1;
tie_graph[891] <= 1'b1;
tie_graph[897] <= 1'b1;
tie_graph[898] <= 1'b1;
tie_graph[900] <= 1'b1;
tie_graph[901] <= 1'b1;
tie_graph[907] <= 1'b1;
tie_graph[908] <= 1'b1;
tie_graph[920] <= 1'b1;
tie_graph[921] <= 1'b1;
tie_graph[926] <= 1'b1;
tie_graph[937] <= 1'b1;
tie_graph[938] <= 1'b1;
tie_graph[943] <= 1'b1;
tie_graph[944] <= 1'b1;
tie_graph[959] <= 1'b1;
tie_graph[960] <= 1'b1;
tie_graph[968] <= 1'b1;
tie_graph[969] <= 1'b1;
tie_graph[974] <= 1'b1;
tie_graph[975] <= 1'b1;
tie_graph[976] <= 1'b1;
tie_graph[980] <= 1'b1;
tie_graph[981] <= 1'b1;
tie_graph[982] <= 1'b1;
tie_graph[987] <= 1'b1;
tie_graph[988] <= 1'b1;
tie_graph[990] <= 1'b1;
tie_graph[991] <= 1'b1;
tie_graph[997] <= 1'b1;
tie_graph[998] <= 1'b1;
tie_graph[1009] <= 1'b1;
tie_graph[1010] <= 1'b1;
tie_graph[1033] <= 1'b1;
tie_graph[1034] <= 1'b1;
tie_graph[1049] <= 1'b1;
tie_graph[1050] <= 1'b1;
tie_graph[1058] <= 1'b1;
tie_graph[1059] <= 1'b1;
tie_graph[1064] <= 1'b1;
tie_graph[1065] <= 1'b1;
tie_graph[1071] <= 1'b1;
tie_graph[1072] <= 1'b1;
tie_graph[1077] <= 1'b1;
tie_graph[1078] <= 1'b1;
tie_graph[1080] <= 1'b1;
tie_graph[1081] <= 1'b1;
tie_graph[1087] <= 1'b1;
tie_graph[1088] <= 1'b1;
tie_graph[1099] <= 1'b1;
tie_graph[1100] <= 1'b1;
tie_graph[1123] <= 1'b1;
tie_graph[1124] <= 1'b1;
tie_graph[1139] <= 1'b1;
tie_graph[1140] <= 1'b1;
tie_graph[1148] <= 1'b1;
tie_graph[1149] <= 1'b1;
tie_graph[1153] <= 1'b1;
tie_graph[1154] <= 1'b1;
tie_graph[1162] <= 1'b1;
tie_graph[1163] <= 1'b1;
tie_graph[1167] <= 1'b1;
tie_graph[1168] <= 1'b1;
tie_graph[1170] <= 1'b1;
tie_graph[1171] <= 1'b1;
tie_graph[1177] <= 1'b1;
tie_graph[1178] <= 1'b1;
tie_graph[1190] <= 1'b1;
tie_graph[1191] <= 1'b1;
tie_graph[1192] <= 1'b1;
tie_graph[1209] <= 1'b1;
tie_graph[1210] <= 1'b1;
tie_graph[1211] <= 1'b1;
tie_graph[1212] <= 1'b1;
tie_graph[1213] <= 1'b1;
tie_graph[1214] <= 1'b1;
tie_graph[1229] <= 1'b1;
tie_graph[1230] <= 1'b1;
tie_graph[1238] <= 1'b1;
tie_graph[1239] <= 1'b1;
tie_graph[1243] <= 1'b1;
tie_graph[1244] <= 1'b1;
tie_graph[1245] <= 1'b1;
tie_graph[1246] <= 1'b1;
tie_graph[1247] <= 1'b1;
tie_graph[1248] <= 1'b1;
tie_graph[1249] <= 1'b1;
tie_graph[1250] <= 1'b1;
tie_graph[1251] <= 1'b1;
tie_graph[1252] <= 1'b1;
tie_graph[1253] <= 1'b1;
tie_graph[1257] <= 1'b1;
tie_graph[1258] <= 1'b1;
tie_graph[1260] <= 1'b1;
tie_graph[1261] <= 1'b1;
tie_graph[1267] <= 1'b1;
tie_graph[1268] <= 1'b1;
tie_graph[1281] <= 1'b1;
tie_graph[1282] <= 1'b1;
tie_graph[1283] <= 1'b1;
tie_graph[1284] <= 1'b1;
tie_graph[1297] <= 1'b1;
tie_graph[1298] <= 1'b1;
tie_graph[1299] <= 1'b1;
tie_graph[1300] <= 1'b1;
tie_graph[1301] <= 1'b1;
tie_graph[1302] <= 1'b1;
tie_graph[1303] <= 1'b1;
tie_graph[1304] <= 1'b1;
tie_graph[1319] <= 1'b1;
tie_graph[1320] <= 1'b1;
tie_graph[1328] <= 1'b1;
tie_graph[1329] <= 1'b1;
tie_graph[1333] <= 1'b1;
tie_graph[1334] <= 1'b1;
tie_graph[1335] <= 1'b1;
tie_graph[1336] <= 1'b1;
tie_graph[1337] <= 1'b1;
tie_graph[1338] <= 1'b1;
tie_graph[1339] <= 1'b1;
tie_graph[1340] <= 1'b1;
tie_graph[1341] <= 1'b1;
tie_graph[1342] <= 1'b1;
tie_graph[1343] <= 1'b1;
tie_graph[1347] <= 1'b1;
tie_graph[1348] <= 1'b1;
tie_graph[1350] <= 1'b1;
tie_graph[1351] <= 1'b1;
tie_graph[1357] <= 1'b1;
tie_graph[1358] <= 1'b1;
tie_graph[1373] <= 1'b1;
tie_graph[1374] <= 1'b1;
tie_graph[1375] <= 1'b1;
tie_graph[1386] <= 1'b1;
tie_graph[1388] <= 1'b1;
tie_graph[1393] <= 1'b1;
tie_graph[1394] <= 1'b1;
tie_graph[1409] <= 1'b1;
tie_graph[1410] <= 1'b1;
tie_graph[1418] <= 1'b1;
tie_graph[1419] <= 1'b1;
tie_graph[1423] <= 1'b1;
tie_graph[1424] <= 1'b1;
tie_graph[1437] <= 1'b1;
tie_graph[1438] <= 1'b1;
tie_graph[1440] <= 1'b1;
tie_graph[1441] <= 1'b1;
tie_graph[1447] <= 1'b1;
tie_graph[1448] <= 1'b1;
tie_graph[1465] <= 1'b1;
tie_graph[1466] <= 1'b1;
tie_graph[1476] <= 1'b1;
tie_graph[1477] <= 1'b1;
tie_graph[1483] <= 1'b1;
tie_graph[1484] <= 1'b1;
tie_graph[1499] <= 1'b1;
tie_graph[1500] <= 1'b1;
tie_graph[1508] <= 1'b1;
tie_graph[1509] <= 1'b1;
tie_graph[1513] <= 1'b1;
tie_graph[1514] <= 1'b1;
tie_graph[1530] <= 1'b1;
tie_graph[1531] <= 1'b1;
tie_graph[1537] <= 1'b1;
tie_graph[1538] <= 1'b1;
tie_graph[1556] <= 1'b1;
tie_graph[1557] <= 1'b1;
tie_graph[1566] <= 1'b1;
tie_graph[1567] <= 1'b1;
tie_graph[1573] <= 1'b1;
tie_graph[1574] <= 1'b1;
tie_graph[1589] <= 1'b1;
tie_graph[1590] <= 1'b1;
tie_graph[1598] <= 1'b1;
tie_graph[1599] <= 1'b1;
tie_graph[1603] <= 1'b1;
tie_graph[1604] <= 1'b1;
tie_graph[1605] <= 1'b1;
tie_graph[1612] <= 1'b1;
tie_graph[1613] <= 1'b1;
tie_graph[1620] <= 1'b1;
tie_graph[1621] <= 1'b1;
tie_graph[1627] <= 1'b1;
tie_graph[1628] <= 1'b1;
tie_graph[1639] <= 1'b1;
tie_graph[1645] <= 1'b1;
tie_graph[1646] <= 1'b1;
tie_graph[1647] <= 1'b1;
tie_graph[1656] <= 1'b1;
tie_graph[1657] <= 1'b1;
tie_graph[1662] <= 1'b1;
tie_graph[1663] <= 1'b1;
tie_graph[1664] <= 1'b1;
tie_graph[1679] <= 1'b1;
tie_graph[1680] <= 1'b1;
tie_graph[1688] <= 1'b1;
tie_graph[1689] <= 1'b1;
tie_graph[1694] <= 1'b1;
tie_graph[1695] <= 1'b1;
tie_graph[1696] <= 1'b1;
tie_graph[1701] <= 1'b1;
tie_graph[1702] <= 1'b1;
tie_graph[1703] <= 1'b1;
tie_graph[1710] <= 1'b1;
tie_graph[1711] <= 1'b1;
tie_graph[1717] <= 1'b1;
tie_graph[1718] <= 1'b1;
tie_graph[1719] <= 1'b1;
tie_graph[1720] <= 1'b1;
tie_graph[1721] <= 1'b1;
tie_graph[1722] <= 1'b1;
tie_graph[1729] <= 1'b1;
tie_graph[1730] <= 1'b1;
tie_graph[1731] <= 1'b1;
tie_graph[1734] <= 1'b1;
tie_graph[1735] <= 1'b1;
tie_graph[1736] <= 1'b1;
tie_graph[1746] <= 1'b1;
tie_graph[1747] <= 1'b1;
tie_graph[1748] <= 1'b1;
tie_graph[1749] <= 1'b1;
tie_graph[1750] <= 1'b1;
tie_graph[1751] <= 1'b1;
tie_graph[1752] <= 1'b1;
tie_graph[1753] <= 1'b1;
tie_graph[1754] <= 1'b1;
tie_graph[1769] <= 1'b1;
tie_graph[1770] <= 1'b1;
tie_graph[1778] <= 1'b1;
tie_graph[1779] <= 1'b1;
tie_graph[1785] <= 1'b1;
tie_graph[1786] <= 1'b1;
tie_graph[1787] <= 1'b1;
tie_graph[1788] <= 1'b1;
tie_graph[1789] <= 1'b1;
tie_graph[1790] <= 1'b1;
tie_graph[1791] <= 1'b1;
tie_graph[1792] <= 1'b1;
tie_graph[1797] <= 1'b1;
tie_graph[1798] <= 1'b1;
tie_graph[1800] <= 1'b1;
tie_graph[1801] <= 1'b1;
tie_graph[1808] <= 1'b1;
tie_graph[1809] <= 1'b1;
tie_graph[1810] <= 1'b1;
tie_graph[1811] <= 1'b1;
tie_graph[1820] <= 1'b1;
tie_graph[1821] <= 1'b1;
tie_graph[1822] <= 1'b1;
tie_graph[1823] <= 1'b1;
tie_graph[1824] <= 1'b1;
tie_graph[1837] <= 1'b1;
tie_graph[1838] <= 1'b1;
tie_graph[1839] <= 1'b1;
tie_graph[1840] <= 1'b1;
tie_graph[1841] <= 1'b1;
tie_graph[1843] <= 1'b1;
tie_graph[1844] <= 1'b1;
tie_graph[1859] <= 1'b1;
tie_graph[1860] <= 1'b1;
tie_graph[1868] <= 1'b1;
tie_graph[1869] <= 1'b1;
tie_graph[1876] <= 1'b1;
tie_graph[1877] <= 1'b1;
tie_graph[1878] <= 1'b1;
tie_graph[1879] <= 1'b1;
tie_graph[1880] <= 1'b1;
tie_graph[1881] <= 1'b1;
tie_graph[1887] <= 1'b1;
tie_graph[1888] <= 1'b1;

				end
			2'b01, 2'b10:
				begin
					win_graph[356] <= 1'b1;
win_graph[357] <= 1'b1;
win_graph[382] <= 1'b1;
win_graph[383] <= 1'b1;
win_graph[392] <= 1'b1;
win_graph[393] <= 1'b1;
win_graph[427] <= 1'b1;
win_graph[428] <= 1'b1;
win_graph[437] <= 1'b1;
win_graph[438] <= 1'b1;
win_graph[447] <= 1'b1;
win_graph[448] <= 1'b1;
win_graph[451] <= 1'b1;
win_graph[452] <= 1'b1;
win_graph[471] <= 1'b1;
win_graph[472] <= 1'b1;
win_graph[478] <= 1'b1;
win_graph[487] <= 1'b1;
win_graph[522] <= 1'b1;
win_graph[523] <= 1'b1;
win_graph[532] <= 1'b1;
win_graph[533] <= 1'b1;
win_graph[542] <= 1'b1;
win_graph[543] <= 1'b1;
win_graph[566] <= 1'b1;
win_graph[567] <= 1'b1;
win_graph[573] <= 1'b1;
win_graph[574] <= 1'b1;
win_graph[581] <= 1'b1;
win_graph[582] <= 1'b1;
win_graph[618] <= 1'b1;
win_graph[619] <= 1'b1;
win_graph[627] <= 1'b1;
win_graph[628] <= 1'b1;
win_graph[636] <= 1'b1;
win_graph[637] <= 1'b1;
win_graph[661] <= 1'b1;
win_graph[662] <= 1'b1;
win_graph[669] <= 1'b1;
win_graph[676] <= 1'b1;
win_graph[713] <= 1'b1;
win_graph[714] <= 1'b1;
win_graph[721] <= 1'b1;
win_graph[722] <= 1'b1;
win_graph[723] <= 1'b1;
win_graph[724] <= 1'b1;
win_graph[731] <= 1'b1;
win_graph[732] <= 1'b1;
win_graph[756] <= 1'b1;
win_graph[757] <= 1'b1;
win_graph[764] <= 1'b1;
win_graph[765] <= 1'b1;
win_graph[770] <= 1'b1;
win_graph[771] <= 1'b1;
win_graph[778] <= 1'b1;
win_graph[779] <= 1'b1;
win_graph[780] <= 1'b1;
win_graph[788] <= 1'b1;
win_graph[789] <= 1'b1;
win_graph[796] <= 1'b1;
win_graph[797] <= 1'b1;
win_graph[808] <= 1'b1;
win_graph[809] <= 1'b1;
win_graph[816] <= 1'b1;
win_graph[817] <= 1'b1;
win_graph[818] <= 1'b1;
win_graph[819] <= 1'b1;
win_graph[826] <= 1'b1;
win_graph[827] <= 1'b1;
win_graph[831] <= 1'b1;
win_graph[832] <= 1'b1;
win_graph[837] <= 1'b1;
win_graph[838] <= 1'b1;
win_graph[841] <= 1'b1;
win_graph[842] <= 1'b1;
win_graph[843] <= 1'b1;
win_graph[851] <= 1'b1;
win_graph[852] <= 1'b1;
win_graph[860] <= 1'b1;
win_graph[865] <= 1'b1;
win_graph[871] <= 1'b1;
win_graph[872] <= 1'b1;
win_graph[873] <= 1'b1;
win_graph[874] <= 1'b1;
win_graph[875] <= 1'b1;
win_graph[876] <= 1'b1;
win_graph[877] <= 1'b1;
win_graph[883] <= 1'b1;
win_graph[884] <= 1'b1;
win_graph[891] <= 1'b1;
win_graph[892] <= 1'b1;
win_graph[904] <= 1'b1;
win_graph[905] <= 1'b1;
win_graph[911] <= 1'b1;
win_graph[914] <= 1'b1;
win_graph[920] <= 1'b1;
win_graph[921] <= 1'b1;
win_graph[926] <= 1'b1;
win_graph[927] <= 1'b1;
win_graph[933] <= 1'b1;
win_graph[935] <= 1'b1;
win_graph[936] <= 1'b1;
win_graph[938] <= 1'b1;
win_graph[939] <= 1'b1;
win_graph[940] <= 1'b1;
win_graph[946] <= 1'b1;
win_graph[947] <= 1'b1;
win_graph[955] <= 1'b1;
win_graph[956] <= 1'b1;
win_graph[959] <= 1'b1;
win_graph[960] <= 1'b1;
win_graph[965] <= 1'b1;
win_graph[966] <= 1'b1;
win_graph[972] <= 1'b1;
win_graph[973] <= 1'b1;
win_graph[978] <= 1'b1;
win_graph[979] <= 1'b1;
win_graph[986] <= 1'b1;
win_graph[987] <= 1'b1;
win_graph[999] <= 1'b1;
win_graph[1000] <= 1'b1;
win_graph[1005] <= 1'b1;
win_graph[1006] <= 1'b1;
win_graph[1009] <= 1'b1;
win_graph[1010] <= 1'b1;
win_graph[1015] <= 1'b1;
win_graph[1016] <= 1'b1;
win_graph[1021] <= 1'b1;
win_graph[1022] <= 1'b1;
win_graph[1028] <= 1'b1;
win_graph[1029] <= 1'b1;
win_graph[1030] <= 1'b1;
win_graph[1034] <= 1'b1;
win_graph[1035] <= 1'b1;
win_graph[1041] <= 1'b1;
win_graph[1042] <= 1'b1;
win_graph[1051] <= 1'b1;
win_graph[1054] <= 1'b1;
win_graph[1059] <= 1'b1;
win_graph[1060] <= 1'b1;
win_graph[1068] <= 1'b1;
win_graph[1069] <= 1'b1;
win_graph[1073] <= 1'b1;
win_graph[1074] <= 1'b1;
win_graph[1081] <= 1'b1;
win_graph[1082] <= 1'b1;
win_graph[1094] <= 1'b1;
win_graph[1095] <= 1'b1;
win_graph[1100] <= 1'b1;
win_graph[1101] <= 1'b1;
win_graph[1104] <= 1'b1;
win_graph[1105] <= 1'b1;
win_graph[1110] <= 1'b1;
win_graph[1111] <= 1'b1;
win_graph[1116] <= 1'b1;
win_graph[1117] <= 1'b1;
win_graph[1123] <= 1'b1;
win_graph[1124] <= 1'b1;
win_graph[1130] <= 1'b1;
win_graph[1131] <= 1'b1;
win_graph[1136] <= 1'b1;
win_graph[1137] <= 1'b1;
win_graph[1146] <= 1'b1;
win_graph[1147] <= 1'b1;
win_graph[1148] <= 1'b1;
win_graph[1149] <= 1'b1;
win_graph[1154] <= 1'b1;
win_graph[1155] <= 1'b1;
win_graph[1163] <= 1'b1;
win_graph[1164] <= 1'b1;
win_graph[1168] <= 1'b1;
win_graph[1169] <= 1'b1;
win_graph[1176] <= 1'b1;
win_graph[1177] <= 1'b1;
win_graph[1190] <= 1'b1;
win_graph[1191] <= 1'b1;
win_graph[1195] <= 1'b1;
win_graph[1200] <= 1'b1;
win_graph[1204] <= 1'b1;
win_graph[1205] <= 1'b1;
win_graph[1211] <= 1'b1;
win_graph[1212] <= 1'b1;
win_graph[1218] <= 1'b1;
win_graph[1225] <= 1'b1;
win_graph[1226] <= 1'b1;
win_graph[1231] <= 1'b1;
win_graph[1232] <= 1'b1;
win_graph[1242] <= 1'b1;
win_graph[1243] <= 1'b1;
win_graph[1248] <= 1'b1;
win_graph[1249] <= 1'b1;
win_graph[1259] <= 1'b1;
win_graph[1260] <= 1'b1;
win_graph[1263] <= 1'b1;
win_graph[1264] <= 1'b1;
win_graph[1271] <= 1'b1;
win_graph[1272] <= 1'b1;
win_graph[1285] <= 1'b1;
win_graph[1286] <= 1'b1;
win_graph[1289] <= 1'b1;
win_graph[1290] <= 1'b1;
win_graph[1295] <= 1'b1;
win_graph[1296] <= 1'b1;
win_graph[1299] <= 1'b1;
win_graph[1300] <= 1'b1;
win_graph[1306] <= 1'b1;
win_graph[1307] <= 1'b1;
win_graph[1312] <= 1'b1;
win_graph[1313] <= 1'b1;
win_graph[1320] <= 1'b1;
win_graph[1321] <= 1'b1;
win_graph[1326] <= 1'b1;
win_graph[1327] <= 1'b1;
win_graph[1337] <= 1'b1;
win_graph[1338] <= 1'b1;
win_graph[1343] <= 1'b1;
win_graph[1344] <= 1'b1;
win_graph[1354] <= 1'b1;
win_graph[1355] <= 1'b1;
win_graph[1358] <= 1'b1;
win_graph[1359] <= 1'b1;
win_graph[1366] <= 1'b1;
win_graph[1367] <= 1'b1;
win_graph[1380] <= 1'b1;
win_graph[1381] <= 1'b1;
win_graph[1384] <= 1'b1;
win_graph[1385] <= 1'b1;
win_graph[1390] <= 1'b1;
win_graph[1391] <= 1'b1;
win_graph[1394] <= 1'b1;
win_graph[1395] <= 1'b1;
win_graph[1401] <= 1'b1;
win_graph[1402] <= 1'b1;
win_graph[1407] <= 1'b1;
win_graph[1408] <= 1'b1;
win_graph[1415] <= 1'b1;
win_graph[1416] <= 1'b1;
win_graph[1421] <= 1'b1;
win_graph[1422] <= 1'b1;
win_graph[1432] <= 1'b1;
win_graph[1433] <= 1'b1;
win_graph[1438] <= 1'b1;
win_graph[1439] <= 1'b1;
win_graph[1449] <= 1'b1;
win_graph[1450] <= 1'b1;
win_graph[1453] <= 1'b1;
win_graph[1454] <= 1'b1;
win_graph[1461] <= 1'b1;
win_graph[1462] <= 1'b1;
win_graph[1475] <= 1'b1;
win_graph[1476] <= 1'b1;
win_graph[1479] <= 1'b1;
win_graph[1480] <= 1'b1;
win_graph[1485] <= 1'b1;
win_graph[1486] <= 1'b1;
win_graph[1489] <= 1'b1;
win_graph[1490] <= 1'b1;
win_graph[1496] <= 1'b1;
win_graph[1497] <= 1'b1;
win_graph[1502] <= 1'b1;
win_graph[1503] <= 1'b1;
win_graph[1510] <= 1'b1;
win_graph[1511] <= 1'b1;
win_graph[1516] <= 1'b1;
win_graph[1517] <= 1'b1;
win_graph[1527] <= 1'b1;
win_graph[1528] <= 1'b1;
win_graph[1534] <= 1'b1;
win_graph[1535] <= 1'b1;
win_graph[1543] <= 1'b1;
win_graph[1544] <= 1'b1;
win_graph[1548] <= 1'b1;
win_graph[1549] <= 1'b1;
win_graph[1556] <= 1'b1;
win_graph[1557] <= 1'b1;
win_graph[1571] <= 1'b1;
win_graph[1572] <= 1'b1;
win_graph[1574] <= 1'b1;
win_graph[1581] <= 1'b1;
win_graph[1583] <= 1'b1;
win_graph[1584] <= 1'b1;
win_graph[1591] <= 1'b1;
win_graph[1592] <= 1'b1;
win_graph[1597] <= 1'b1;
win_graph[1598] <= 1'b1;
win_graph[1605] <= 1'b1;
win_graph[1606] <= 1'b1;
win_graph[1622] <= 1'b1;
win_graph[1623] <= 1'b1;
win_graph[1629] <= 1'b1;
win_graph[1630] <= 1'b1;
win_graph[1638] <= 1'b1;
win_graph[1639] <= 1'b1;
win_graph[1643] <= 1'b1;
win_graph[1644] <= 1'b1;
win_graph[1651] <= 1'b1;
win_graph[1652] <= 1'b1;
win_graph[1666] <= 1'b1;
win_graph[1667] <= 1'b1;
win_graph[1668] <= 1'b1;
win_graph[1669] <= 1'b1;
win_graph[1676] <= 1'b1;
win_graph[1677] <= 1'b1;
win_graph[1678] <= 1'b1;
win_graph[1679] <= 1'b1;
win_graph[1686] <= 1'b1;
win_graph[1687] <= 1'b1;
win_graph[1692] <= 1'b1;
win_graph[1693] <= 1'b1;
win_graph[1700] <= 1'b1;
win_graph[1701] <= 1'b1;
win_graph[1717] <= 1'b1;
win_graph[1718] <= 1'b1;
win_graph[1725] <= 1'b1;
win_graph[1726] <= 1'b1;
win_graph[1732] <= 1'b1;
win_graph[1733] <= 1'b1;
win_graph[1738] <= 1'b1;
win_graph[1739] <= 1'b1;
win_graph[1740] <= 1'b1;
win_graph[1745] <= 1'b1;
win_graph[1746] <= 1'b1;
win_graph[1747] <= 1'b1;
win_graph[1761] <= 1'b1;
win_graph[1762] <= 1'b1;
win_graph[1763] <= 1'b1;
win_graph[1764] <= 1'b1;
win_graph[1771] <= 1'b1;
win_graph[1772] <= 1'b1;
win_graph[1773] <= 1'b1;
win_graph[1774] <= 1'b1;
win_graph[1781] <= 1'b1;
win_graph[1782] <= 1'b1;
win_graph[1787] <= 1'b1;
win_graph[1788] <= 1'b1;
win_graph[1795] <= 1'b1;
win_graph[1796] <= 1'b1;
win_graph[1812] <= 1'b1;
win_graph[1813] <= 1'b1;
win_graph[1821] <= 1'b1;
win_graph[1822] <= 1'b1;
win_graph[1823] <= 1'b1;
win_graph[1824] <= 1'b1;
win_graph[1825] <= 1'b1;
win_graph[1826] <= 1'b1;
win_graph[1827] <= 1'b1;
win_graph[1834] <= 1'b1;
win_graph[1835] <= 1'b1;
win_graph[1836] <= 1'b1;
win_graph[1837] <= 1'b1;
win_graph[1838] <= 1'b1;
win_graph[1839] <= 1'b1;
win_graph[1840] <= 1'b1;
win_graph[1841] <= 1'b1;
win_graph[1842] <= 1'b1;
win_graph[1857] <= 1'b1;
win_graph[1858] <= 1'b1;
win_graph[1867] <= 1'b1;
win_graph[1868] <= 1'b1;
win_graph[1876] <= 1'b1;
win_graph[1877] <= 1'b1;
win_graph[1882] <= 1'b1;
win_graph[1883] <= 1'b1;
win_graph[1890] <= 1'b1;
win_graph[1891] <= 1'b1;
win_graph[1896] <= 1'b1;
win_graph[1897] <= 1'b1;
win_graph[1907] <= 1'b1;
win_graph[1908] <= 1'b1;
win_graph[1918] <= 1'b1;
win_graph[1919] <= 1'b1;
win_graph[1920] <= 1'b1;
win_graph[1930] <= 1'b1;
win_graph[1931] <= 1'b1;
win_graph[1932] <= 1'b1;
win_graph[1933] <= 1'b1;
win_graph[1934] <= 1'b1;
win_graph[1936] <= 1'b1;
win_graph[1937] <= 1'b1;
win_graph[1952] <= 1'b1;
win_graph[1953] <= 1'b1;
win_graph[1962] <= 1'b1;
win_graph[1963] <= 1'b1;
win_graph[1971] <= 1'b1;
win_graph[1972] <= 1'b1;
win_graph[1978] <= 1'b1;
win_graph[1985] <= 1'b1;
win_graph[1986] <= 1'b1;
win_graph[1991] <= 1'b1;
win_graph[1992] <= 1'b1;

				end
	 
	 endcase
end
else
		begin

		tie_graph <= 1'b0;
		win_graph <= 1'b0;
		end
end
endmodule