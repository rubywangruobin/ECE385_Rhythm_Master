module dropper_thirty_nine39(input Reset, frame_clk, 
						 input logic [7:0] keycode,keycode_second,
						 output [9:0] drop39X, drop39Y,
						 output [1599:0] arrow39,
						 output logic score39);
	logic [9:0] arrow_X_Pos, arrow_Y_Pos, arrow_Y_Motion;
	logic [11:0] counter;
    parameter [9:0] X_start=500;  // Center position on the X axis
    parameter [9:0] Y_start=100;  // Center position on the Y axis
    parameter [9:0] Y_Max=400;     // Bottommost point on the Y axis
	 logic finish_on;
	 enum logic [3:0] {Halted, Normal, End} State, Next_state;
	 
	 always_ff @ (posedge frame_clk )
    begin
		if(Reset)
		begin
			State <= Halted;
		end	
		else if(State == Halted)
		begin
			counter = 0;
			score39 = 0;
			arrow_Y_Motion = 0; 
			arrow_Y_Pos = Y_start;
			State <= Next_state;
		end
		else if(State == Normal)
			begin
				if(counter <2800)
					counter = counter + 1;
				else
					begin
						arrow_Y_Motion = 1;
						if ((arrow_Y_Pos + 40) >= Y_Max)
							score39 = 1'b0;	
						else if ((keycode == 8'h4f|| keycode_second == 8'h4f) & (arrow_Y_Pos + 40 >= 340) & (arrow_Y_Pos + 40 < 400))
							score39 = 1'b1;
						else
						begin
							arrow_Y_Pos = (arrow_Y_Pos + arrow_Y_Motion); 
							counter = counter + 1;
						end
					end
				State <= Next_state;
			end
		else
			State <= Next_state;
    end
	 
	 always_comb
	 begin
		Next_state = State;
		finish_on = 1'b0;
		arrow_X_Pos = X_start;
		unique case(State)
			Halted:
			begin
				finish_on = 1'b0;
				if(keycode == 8'h2c)
					Next_state = Normal;
			end
			Normal:
				begin
				if(counter < 2800)
				begin
					Next_state = Normal;
					end
				else
					begin
						if ( (arrow_Y_Pos + 40) >= Y_Max )  
							begin
									finish_on = 1'b1; 
									Next_state = End;
							end
						 else if ((keycode == 8'h4f|| keycode_second == 8'h4f) & (arrow_Y_Pos + 40 >= 340) & (arrow_Y_Pos + 40 < 400))
							begin
									finish_on = 1'b1;
									Next_state = End;
							end
						 else
							begin
								  Next_state = Normal;
							end
					end
				end
			End:
				begin
				finish_on = 1;
				if(keycode == 8'h01)
					Next_state = Halted;
				end
		endcase
					
	 end
    assign drop39X = arrow_X_Pos;
   
    assign drop39Y = arrow_Y_Pos;
	 always_comb
	 begin
	 arrow39 <= 1'b0;
	 if(finish_on == 0)
	 begin
	 arrow39[420] <= 1'b1;
arrow39[421] <= 1'b1;
arrow39[460] <= 1'b1;
arrow39[461] <= 1'b1;
arrow39[500] <= 1'b1;
arrow39[501] <= 1'b1;
arrow39[502] <= 1'b1;
arrow39[503] <= 1'b1;
arrow39[540] <= 1'b1;
arrow39[541] <= 1'b1;
arrow39[542] <= 1'b1;
arrow39[543] <= 1'b1;
arrow39[580] <= 1'b1;
arrow39[581] <= 1'b1;
arrow39[582] <= 1'b1;
arrow39[583] <= 1'b1;
arrow39[584] <= 1'b1;
arrow39[585] <= 1'b1;
arrow39[620] <= 1'b1;
arrow39[621] <= 1'b1;
arrow39[622] <= 1'b1;
arrow39[623] <= 1'b1;
arrow39[624] <= 1'b1;
arrow39[625] <= 1'b1;
arrow39[648] <= 1'b1;
arrow39[649] <= 1'b1;
arrow39[650] <= 1'b1;
arrow39[651] <= 1'b1;
arrow39[652] <= 1'b1;
arrow39[653] <= 1'b1;
arrow39[654] <= 1'b1;
arrow39[655] <= 1'b1;
arrow39[656] <= 1'b1;
arrow39[657] <= 1'b1;
arrow39[658] <= 1'b1;
arrow39[659] <= 1'b1;
arrow39[660] <= 1'b1;
arrow39[661] <= 1'b1;
arrow39[662] <= 1'b1;
arrow39[663] <= 1'b1;
arrow39[664] <= 1'b1;
arrow39[665] <= 1'b1;
arrow39[666] <= 1'b1;
arrow39[667] <= 1'b1;
arrow39[688] <= 1'b1;
arrow39[689] <= 1'b1;
arrow39[690] <= 1'b1;
arrow39[691] <= 1'b1;
arrow39[692] <= 1'b1;
arrow39[693] <= 1'b1;
arrow39[694] <= 1'b1;
arrow39[695] <= 1'b1;
arrow39[696] <= 1'b1;
arrow39[697] <= 1'b1;
arrow39[698] <= 1'b1;
arrow39[699] <= 1'b1;
arrow39[700] <= 1'b1;
arrow39[701] <= 1'b1;
arrow39[702] <= 1'b1;
arrow39[703] <= 1'b1;
arrow39[704] <= 1'b1;
arrow39[705] <= 1'b1;
arrow39[706] <= 1'b1;
arrow39[707] <= 1'b1;
arrow39[728] <= 1'b1;
arrow39[729] <= 1'b1;
arrow39[730] <= 1'b1;
arrow39[731] <= 1'b1;
arrow39[732] <= 1'b1;
arrow39[733] <= 1'b1;
arrow39[734] <= 1'b1;
arrow39[735] <= 1'b1;
arrow39[736] <= 1'b1;
arrow39[737] <= 1'b1;
arrow39[738] <= 1'b1;
arrow39[739] <= 1'b1;
arrow39[740] <= 1'b1;
arrow39[741] <= 1'b1;
arrow39[742] <= 1'b1;
arrow39[743] <= 1'b1;
arrow39[744] <= 1'b1;
arrow39[745] <= 1'b1;
arrow39[746] <= 1'b1;
arrow39[747] <= 1'b1;
arrow39[748] <= 1'b1;
arrow39[749] <= 1'b1;
arrow39[768] <= 1'b1;
arrow39[769] <= 1'b1;
arrow39[770] <= 1'b1;
arrow39[771] <= 1'b1;
arrow39[772] <= 1'b1;
arrow39[773] <= 1'b1;
arrow39[774] <= 1'b1;
arrow39[775] <= 1'b1;
arrow39[776] <= 1'b1;
arrow39[777] <= 1'b1;
arrow39[778] <= 1'b1;
arrow39[779] <= 1'b1;
arrow39[780] <= 1'b1;
arrow39[781] <= 1'b1;
arrow39[782] <= 1'b1;
arrow39[783] <= 1'b1;
arrow39[784] <= 1'b1;
arrow39[785] <= 1'b1;
arrow39[786] <= 1'b1;
arrow39[787] <= 1'b1;
arrow39[788] <= 1'b1;
arrow39[789] <= 1'b1;
arrow39[808] <= 1'b1;
arrow39[809] <= 1'b1;
arrow39[810] <= 1'b1;
arrow39[811] <= 1'b1;
arrow39[812] <= 1'b1;
arrow39[813] <= 1'b1;
arrow39[814] <= 1'b1;
arrow39[815] <= 1'b1;
arrow39[816] <= 1'b1;
arrow39[817] <= 1'b1;
arrow39[818] <= 1'b1;
arrow39[819] <= 1'b1;
arrow39[820] <= 1'b1;
arrow39[821] <= 1'b1;
arrow39[822] <= 1'b1;
arrow39[823] <= 1'b1;
arrow39[824] <= 1'b1;
arrow39[825] <= 1'b1;
arrow39[826] <= 1'b1;
arrow39[827] <= 1'b1;
arrow39[848] <= 1'b1;
arrow39[849] <= 1'b1;
arrow39[850] <= 1'b1;
arrow39[851] <= 1'b1;
arrow39[852] <= 1'b1;
arrow39[853] <= 1'b1;
arrow39[854] <= 1'b1;
arrow39[855] <= 1'b1;
arrow39[856] <= 1'b1;
arrow39[857] <= 1'b1;
arrow39[858] <= 1'b1;
arrow39[859] <= 1'b1;
arrow39[860] <= 1'b1;
arrow39[861] <= 1'b1;
arrow39[862] <= 1'b1;
arrow39[863] <= 1'b1;
arrow39[864] <= 1'b1;
arrow39[865] <= 1'b1;
arrow39[866] <= 1'b1;
arrow39[867] <= 1'b1;
arrow39[900] <= 1'b1;
arrow39[901] <= 1'b1;
arrow39[902] <= 1'b1;
arrow39[903] <= 1'b1;
arrow39[904] <= 1'b1;
arrow39[905] <= 1'b1;
arrow39[940] <= 1'b1;
arrow39[941] <= 1'b1;
arrow39[942] <= 1'b1;
arrow39[943] <= 1'b1;
arrow39[944] <= 1'b1;
arrow39[945] <= 1'b1;
arrow39[980] <= 1'b1;
arrow39[981] <= 1'b1;
arrow39[982] <= 1'b1;
arrow39[983] <= 1'b1;
arrow39[1020] <= 1'b1;
arrow39[1021] <= 1'b1;
arrow39[1022] <= 1'b1;
arrow39[1023] <= 1'b1;
arrow39[1060] <= 1'b1;
arrow39[1061] <= 1'b1;
arrow39[1100] <= 1'b1;
arrow39[1101] <= 1'b1;


	 end
   else
		 arrow39 <= 1'b0;
end
endmodule