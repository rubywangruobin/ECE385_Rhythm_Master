module palette(input address, output logic[23:0] RGB);
always_comb begin
			case (address)
			
endcase
end
endmodule
