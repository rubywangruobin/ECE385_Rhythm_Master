module pika (input Reset, frame_clk, 
				 input logic [7:0] keycode,
				 output [17249:0] pika_color);
				 
				 
				 
	enum logic [7:0] {Start_state, Halted, move1, move2, move3, move4, move5,
							move6, move7, move8, move9, move10, move11,
							move12, move13, move14, move15, move16, move17, move18,
							move19, move20, move21, move22, move23, move24, move25,
							move26, move27, move28, move29, move30, move31, move32,
							move33, move34, move35, move36, move37, move38, move39,
							move40, move41, move42, move43, move44, move45, move46, 
							move47, move48, move49, move50, move51, move52, move53,
							move54, move55, move56, move57, move58, move59, move60,
							move61, move62, move63, move64, move65, move66, move67,
							move68, move69, move70, move71, move72, move73, move74,
							move75, move76, move77, move78, move79} State, Next_state;
	always_ff @ (posedge frame_clk) begin
		if(Reset)
			State <= Start_state;
		else
			State <= Next_state;
	end
	
	always_comb
	begin
	Next_state = State;
	pika_color = 0;
	unique case (State)
		Start_state:
			if(keycode == 8'h2c)
			  Next_state = Halted;
		Halted:
			Next_state = move1;
		move1:
			Next_state = move2;
		move2:
			Next_state = move3;
		move3:
			Next_state = move4;
		move4:
			Next_state = move5;
		move5:
			Next_state = move6;
		move6:
			Next_state = move7;
		move7:
			Next_state = move8;
		move8:
			Next_state = move9;
		move9:
			Next_state = move10;
		move10:
			Next_state = move11;
		
	  move11:
		Next_state = move12;
	  move12:
		Next_state = move13;
	  move13:
		Next_state = move14;
	  move14:
		Next_state = move15;
	  move15:
		Next_state = move16;
	  move16:
		Next_state = move17;
	  move17:
		Next_state = move18;
	  move18:
		Next_state = move19;
	  move19:
		Next_state = move20;
	  move20:
		Next_state = move21;
	  move21:
		Next_state = move22;
	  move22:
		Next_state = move23;
	  move23:
		Next_state = move24;
	  move24:
		Next_state = move25;
	  move25:
		Next_state = move26;
	  move26:
		Next_state = move27;
	  move27:
		Next_state = move28;
	  move28:
		Next_state = move29;
	  move29:
		Next_state = move30;
	  move30:
		Next_state = move31;
	  move31:
		Next_state = move32;
	  move32:
		Next_state = move33;
	  move33:
		Next_state = move34;
	  move34:
		Next_state = move35;
	  move35:
		Next_state = move36;
	  move36:
		Next_state = move37;
	  move37:
		Next_state = move38;
	  move38:
		Next_state = move39;
	  move39:
		Next_state = move40;
	  move40:
		Next_state = move41;
	  move41:
		Next_state = move42;
	  move42:
		Next_state = move43;
	  move43:
		Next_state = move44;
	  move44:
		Next_state = move45;
	  move45:
		Next_state = move46;
	  move46:
		Next_state = move47;
	  move47:
		Next_state = move48;
	  move48:
		Next_state = move49;
	  move49:
		Next_state = move50;
	  move50:
		Next_state = move51;
	  move51:
		Next_state = move52;
	  move52:
		Next_state = move53;
	  move53:
		Next_state = move54;
	  move54:
		Next_state = move55;
	  move55:
		Next_state = move56;
	  move56:
		Next_state = move57;
	  move57:
		Next_state = move58;
	  move58:
		Next_state = move59;
	  move59:
		Next_state = move60;
	  move60:
		Next_state = move61;
	  move61:
		Next_state = move62;
	  move62:
		Next_state = move63;
	  move63:
		Next_state = move64;
	  move64:
		Next_state = move65;
	  move65:
		Next_state = move66;
	  move66:
		Next_state = move67;
	  move67:
		Next_state = move68;
	  move68:
		Next_state = move69;
	  move69:
		Next_state = move70;
	  move70:
		Next_state = move71;
	  move71:
		Next_state = move72;
	  move72:
		Next_state = move73;
	  move73:
		Next_state = move74;
	  move74:
		Next_state = move75;
	  move75:
		Next_state = move76;
	  move76:
		Next_state = move77;
	  move77:
		Next_state = move78;
	  move78:
		Next_state = move79;
	  move79:
		Next_state = Halted;
	  
		default:;
		
	endcase
	case(State)
		Start_state, Halted, move1, move2, move3, move4, move5, move6, move7, move8, move9:
		begin
			pika_color[943] <= 1'b1;
pika_color[944] <= 1'b1;
pika_color[945] <= 1'b1;
pika_color[946] <= 1'b1;
pika_color[1058] <= 1'b1;
pika_color[1059] <= 1'b1;
pika_color[1060] <= 1'b1;
pika_color[1061] <= 1'b1;
pika_color[1062] <= 1'b1;
pika_color[1172] <= 1'b1;
pika_color[1173] <= 1'b1;
pika_color[1174] <= 1'b1;
pika_color[1175] <= 1'b1;
pika_color[1176] <= 1'b1;
pika_color[1177] <= 1'b1;
pika_color[1178] <= 1'b1;
pika_color[1274] <= 1'b1;
pika_color[1275] <= 1'b1;
pika_color[1276] <= 1'b1;
pika_color[1287] <= 1'b1;
pika_color[1288] <= 1'b1;
pika_color[1289] <= 1'b1;
pika_color[1290] <= 1'b1;
pika_color[1291] <= 1'b1;
pika_color[1292] <= 1'b1;
pika_color[1293] <= 1'b1;
pika_color[1294] <= 1'b1;
pika_color[1295] <= 1'b1;
pika_color[1389] <= 1'b1;
pika_color[1391] <= 1'b1;
pika_color[1392] <= 1'b1;
pika_color[1402] <= 1'b1;
pika_color[1403] <= 1'b1;
pika_color[1404] <= 1'b1;
pika_color[1405] <= 1'b1;
pika_color[1406] <= 1'b1;
pika_color[1407] <= 1'b1;
pika_color[1408] <= 1'b1;
pika_color[1409] <= 1'b1;
pika_color[1410] <= 1'b1;
pika_color[1411] <= 1'b1;
pika_color[1504] <= 1'b1;
pika_color[1507] <= 1'b1;
pika_color[1508] <= 1'b1;
pika_color[1518] <= 1'b1;
pika_color[1519] <= 1'b1;
pika_color[1520] <= 1'b1;
pika_color[1521] <= 1'b1;
pika_color[1522] <= 1'b1;
pika_color[1523] <= 1'b1;
pika_color[1524] <= 1'b1;
pika_color[1526] <= 1'b1;
pika_color[1527] <= 1'b1;
pika_color[1619] <= 1'b1;
pika_color[1623] <= 1'b1;
pika_color[1624] <= 1'b1;
pika_color[1633] <= 1'b1;
pika_color[1634] <= 1'b1;
pika_color[1635] <= 1'b1;
pika_color[1636] <= 1'b1;
pika_color[1637] <= 1'b1;
pika_color[1638] <= 1'b1;
pika_color[1639] <= 1'b1;
pika_color[1643] <= 1'b1;
pika_color[1734] <= 1'b1;
pika_color[1739] <= 1'b1;
pika_color[1740] <= 1'b1;
pika_color[1748] <= 1'b1;
pika_color[1749] <= 1'b1;
pika_color[1750] <= 1'b1;
pika_color[1751] <= 1'b1;
pika_color[1752] <= 1'b1;
pika_color[1753] <= 1'b1;
pika_color[1754] <= 1'b1;
pika_color[1759] <= 1'b1;
pika_color[1849] <= 1'b1;
pika_color[1855] <= 1'b1;
pika_color[1856] <= 1'b1;
pika_color[1864] <= 1'b1;
pika_color[1865] <= 1'b1;
pika_color[1866] <= 1'b1;
pika_color[1867] <= 1'b1;
pika_color[1868] <= 1'b1;
pika_color[1869] <= 1'b1;
pika_color[1874] <= 1'b1;
pika_color[1875] <= 1'b1;
pika_color[1964] <= 1'b1;
pika_color[1971] <= 1'b1;
pika_color[1972] <= 1'b1;
pika_color[1979] <= 1'b1;
pika_color[1980] <= 1'b1;
pika_color[1981] <= 1'b1;
pika_color[1982] <= 1'b1;
pika_color[1983] <= 1'b1;
pika_color[1984] <= 1'b1;
pika_color[1990] <= 1'b1;
pika_color[1991] <= 1'b1;
pika_color[2079] <= 1'b1;
pika_color[2087] <= 1'b1;
pika_color[2088] <= 1'b1;
pika_color[2095] <= 1'b1;
pika_color[2096] <= 1'b1;
pika_color[2097] <= 1'b1;
pika_color[2098] <= 1'b1;
pika_color[2106] <= 1'b1;
pika_color[2107] <= 1'b1;
pika_color[2194] <= 1'b1;
pika_color[2203] <= 1'b1;
pika_color[2204] <= 1'b1;
pika_color[2210] <= 1'b1;
pika_color[2211] <= 1'b1;
pika_color[2212] <= 1'b1;
pika_color[2213] <= 1'b1;
pika_color[2223] <= 1'b1;
pika_color[2309] <= 1'b1;
pika_color[2320] <= 1'b1;
pika_color[2325] <= 1'b1;
pika_color[2326] <= 1'b1;
pika_color[2327] <= 1'b1;
pika_color[2328] <= 1'b1;
pika_color[2338] <= 1'b1;
pika_color[2339] <= 1'b1;
pika_color[2424] <= 1'b1;
pika_color[2435] <= 1'b1;
pika_color[2436] <= 1'b1;
pika_color[2440] <= 1'b1;
pika_color[2441] <= 1'b1;
pika_color[2442] <= 1'b1;
pika_color[2443] <= 1'b1;
pika_color[2454] <= 1'b1;
pika_color[2539] <= 1'b1;
pika_color[2551] <= 1'b1;
pika_color[2552] <= 1'b1;
pika_color[2556] <= 1'b1;
pika_color[2557] <= 1'b1;
pika_color[2558] <= 1'b1;
pika_color[2569] <= 1'b1;
pika_color[2570] <= 1'b1;
pika_color[2654] <= 1'b1;
pika_color[2667] <= 1'b1;
pika_color[2671] <= 1'b1;
pika_color[2672] <= 1'b1;
pika_color[2673] <= 1'b1;
pika_color[2685] <= 1'b1;
pika_color[2769] <= 1'b1;
pika_color[2783] <= 1'b1;
pika_color[2787] <= 1'b1;
pika_color[2788] <= 1'b1;
pika_color[2801] <= 1'b1;
pika_color[2884] <= 1'b1;
pika_color[2898] <= 1'b1;
pika_color[2899] <= 1'b1;
pika_color[2902] <= 1'b1;
pika_color[2903] <= 1'b1;
pika_color[2916] <= 1'b1;
pika_color[2917] <= 1'b1;
pika_color[2999] <= 1'b1;
pika_color[3000] <= 1'b1;
pika_color[3014] <= 1'b1;
pika_color[3018] <= 1'b1;
pika_color[3032] <= 1'b1;
pika_color[3115] <= 1'b1;
pika_color[3129] <= 1'b1;
pika_color[3130] <= 1'b1;
pika_color[3133] <= 1'b1;
pika_color[3148] <= 1'b1;
pika_color[3230] <= 1'b1;
pika_color[3245] <= 1'b1;
pika_color[3246] <= 1'b1;
pika_color[3249] <= 1'b1;
pika_color[3263] <= 1'b1;
pika_color[3345] <= 1'b1;
pika_color[3361] <= 1'b1;
pika_color[3362] <= 1'b1;
pika_color[3364] <= 1'b1;
pika_color[3365] <= 1'b1;
pika_color[3378] <= 1'b1;
pika_color[3379] <= 1'b1;
pika_color[3460] <= 1'b1;
pika_color[3477] <= 1'b1;
pika_color[3478] <= 1'b1;
pika_color[3480] <= 1'b1;
pika_color[3494] <= 1'b1;
pika_color[3575] <= 1'b1;
pika_color[3593] <= 1'b1;
pika_color[3595] <= 1'b1;
pika_color[3596] <= 1'b1;
pika_color[3609] <= 1'b1;
pika_color[3610] <= 1'b1;
pika_color[3690] <= 1'b1;
pika_color[3691] <= 1'b1;
pika_color[3708] <= 1'b1;
pika_color[3709] <= 1'b1;
pika_color[3711] <= 1'b1;
pika_color[3712] <= 1'b1;
pika_color[3725] <= 1'b1;
pika_color[3806] <= 1'b1;
pika_color[3824] <= 1'b1;
pika_color[3825] <= 1'b1;
pika_color[3827] <= 1'b1;
pika_color[3840] <= 1'b1;
pika_color[3841] <= 1'b1;
pika_color[3921] <= 1'b1;
pika_color[3940] <= 1'b1;
pika_color[3942] <= 1'b1;
pika_color[3943] <= 1'b1;
pika_color[3956] <= 1'b1;
pika_color[4036] <= 1'b1;
pika_color[4055] <= 1'b1;
pika_color[4056] <= 1'b1;
pika_color[4058] <= 1'b1;
pika_color[4059] <= 1'b1;
pika_color[4071] <= 1'b1;
pika_color[4151] <= 1'b1;
pika_color[4171] <= 1'b1;
pika_color[4174] <= 1'b1;
pika_color[4187] <= 1'b1;
pika_color[4266] <= 1'b1;
pika_color[4286] <= 1'b1;
pika_color[4287] <= 1'b1;
pika_color[4289] <= 1'b1;
pika_color[4302] <= 1'b1;
pika_color[4309] <= 1'b1;
pika_color[4310] <= 1'b1;
pika_color[4311] <= 1'b1;
pika_color[4312] <= 1'b1;
pika_color[4313] <= 1'b1;
pika_color[4381] <= 1'b1;
pika_color[4402] <= 1'b1;
pika_color[4404] <= 1'b1;
pika_color[4405] <= 1'b1;
pika_color[4417] <= 1'b1;
pika_color[4418] <= 1'b1;
pika_color[4419] <= 1'b1;
pika_color[4420] <= 1'b1;
pika_color[4421] <= 1'b1;
pika_color[4422] <= 1'b1;
pika_color[4423] <= 1'b1;
pika_color[4428] <= 1'b1;
pika_color[4429] <= 1'b1;
pika_color[4430] <= 1'b1;
pika_color[4431] <= 1'b1;
pika_color[4432] <= 1'b1;
pika_color[4433] <= 1'b1;
pika_color[4434] <= 1'b1;
pika_color[4462] <= 1'b1;
pika_color[4463] <= 1'b1;
pika_color[4464] <= 1'b1;
pika_color[4465] <= 1'b1;
pika_color[4466] <= 1'b1;
pika_color[4467] <= 1'b1;
pika_color[4468] <= 1'b1;
pika_color[4469] <= 1'b1;
pika_color[4470] <= 1'b1;
pika_color[4471] <= 1'b1;
pika_color[4472] <= 1'b1;
pika_color[4473] <= 1'b1;
pika_color[4474] <= 1'b1;
pika_color[4496] <= 1'b1;
pika_color[4497] <= 1'b1;
pika_color[4517] <= 1'b1;
pika_color[4518] <= 1'b1;
pika_color[4520] <= 1'b1;
pika_color[4521] <= 1'b1;
pika_color[4533] <= 1'b1;
pika_color[4549] <= 1'b1;
pika_color[4550] <= 1'b1;
pika_color[4551] <= 1'b1;
pika_color[4552] <= 1'b1;
pika_color[4553] <= 1'b1;
pika_color[4573] <= 1'b1;
pika_color[4574] <= 1'b1;
pika_color[4575] <= 1'b1;
pika_color[4576] <= 1'b1;
pika_color[4577] <= 1'b1;
pika_color[4588] <= 1'b1;
pika_color[4589] <= 1'b1;
pika_color[4590] <= 1'b1;
pika_color[4591] <= 1'b1;
pika_color[4592] <= 1'b1;
pika_color[4593] <= 1'b1;
pika_color[4612] <= 1'b1;
pika_color[4633] <= 1'b1;
pika_color[4634] <= 1'b1;
pika_color[4636] <= 1'b1;
pika_color[4668] <= 1'b1;
pika_color[4669] <= 1'b1;
pika_color[4687] <= 1'b1;
pika_color[4688] <= 1'b1;
pika_color[4708] <= 1'b1;
pika_color[4709] <= 1'b1;
pika_color[4710] <= 1'b1;
pika_color[4711] <= 1'b1;
pika_color[4712] <= 1'b1;
pika_color[4727] <= 1'b1;
pika_color[4749] <= 1'b1;
pika_color[4752] <= 1'b1;
pika_color[4785] <= 1'b1;
pika_color[4786] <= 1'b1;
pika_color[4787] <= 1'b1;
pika_color[4800] <= 1'b1;
pika_color[4801] <= 1'b1;
pika_color[4822] <= 1'b1;
pika_color[4823] <= 1'b1;
pika_color[4824] <= 1'b1;
pika_color[4825] <= 1'b1;
pika_color[4826] <= 1'b1;
pika_color[4827] <= 1'b1;
pika_color[4828] <= 1'b1;
pika_color[4829] <= 1'b1;
pika_color[4842] <= 1'b1;
pika_color[4864] <= 1'b1;
pika_color[4865] <= 1'b1;
pika_color[4867] <= 1'b1;
pika_color[4902] <= 1'b1;
pika_color[4903] <= 1'b1;
pika_color[4912] <= 1'b1;
pika_color[4913] <= 1'b1;
pika_color[4914] <= 1'b1;
pika_color[4915] <= 1'b1;
pika_color[4936] <= 1'b1;
pika_color[4937] <= 1'b1;
pika_color[4938] <= 1'b1;
pika_color[4939] <= 1'b1;
pika_color[4940] <= 1'b1;
pika_color[4941] <= 1'b1;
pika_color[4942] <= 1'b1;
pika_color[4943] <= 1'b1;
pika_color[4944] <= 1'b1;
pika_color[4957] <= 1'b1;
pika_color[4980] <= 1'b1;
pika_color[4981] <= 1'b1;
pika_color[4983] <= 1'b1;
pika_color[5019] <= 1'b1;
pika_color[5020] <= 1'b1;
pika_color[5022] <= 1'b1;
pika_color[5023] <= 1'b1;
pika_color[5024] <= 1'b1;
pika_color[5025] <= 1'b1;
pika_color[5026] <= 1'b1;
pika_color[5027] <= 1'b1;
pika_color[5050] <= 1'b1;
pika_color[5051] <= 1'b1;
pika_color[5052] <= 1'b1;
pika_color[5053] <= 1'b1;
pika_color[5054] <= 1'b1;
pika_color[5055] <= 1'b1;
pika_color[5056] <= 1'b1;
pika_color[5057] <= 1'b1;
pika_color[5058] <= 1'b1;
pika_color[5059] <= 1'b1;
pika_color[5073] <= 1'b1;
pika_color[5096] <= 1'b1;
pika_color[5097] <= 1'b1;
pika_color[5098] <= 1'b1;
pika_color[5099] <= 1'b1;
pika_color[5135] <= 1'b1;
pika_color[5136] <= 1'b1;
pika_color[5137] <= 1'b1;
pika_color[5164] <= 1'b1;
pika_color[5165] <= 1'b1;
pika_color[5166] <= 1'b1;
pika_color[5167] <= 1'b1;
pika_color[5168] <= 1'b1;
pika_color[5169] <= 1'b1;
pika_color[5170] <= 1'b1;
pika_color[5171] <= 1'b1;
pika_color[5172] <= 1'b1;
pika_color[5173] <= 1'b1;
pika_color[5174] <= 1'b1;
pika_color[5188] <= 1'b1;
pika_color[5212] <= 1'b1;
pika_color[5213] <= 1'b1;
pika_color[5278] <= 1'b1;
pika_color[5279] <= 1'b1;
pika_color[5280] <= 1'b1;
pika_color[5281] <= 1'b1;
pika_color[5282] <= 1'b1;
pika_color[5283] <= 1'b1;
pika_color[5284] <= 1'b1;
pika_color[5285] <= 1'b1;
pika_color[5286] <= 1'b1;
pika_color[5287] <= 1'b1;
pika_color[5288] <= 1'b1;
pika_color[5303] <= 1'b1;
pika_color[5304] <= 1'b1;
pika_color[5326] <= 1'b1;
pika_color[5327] <= 1'b1;
pika_color[5393] <= 1'b1;
pika_color[5394] <= 1'b1;
pika_color[5395] <= 1'b1;
pika_color[5396] <= 1'b1;
pika_color[5397] <= 1'b1;
pika_color[5398] <= 1'b1;
pika_color[5399] <= 1'b1;
pika_color[5400] <= 1'b1;
pika_color[5401] <= 1'b1;
pika_color[5420] <= 1'b1;
pika_color[5421] <= 1'b1;
pika_color[5441] <= 1'b1;
pika_color[5507] <= 1'b1;
pika_color[5508] <= 1'b1;
pika_color[5509] <= 1'b1;
pika_color[5510] <= 1'b1;
pika_color[5511] <= 1'b1;
pika_color[5512] <= 1'b1;
pika_color[5513] <= 1'b1;
pika_color[5514] <= 1'b1;
pika_color[5515] <= 1'b1;
pika_color[5536] <= 1'b1;
pika_color[5556] <= 1'b1;
pika_color[5621] <= 1'b1;
pika_color[5622] <= 1'b1;
pika_color[5623] <= 1'b1;
pika_color[5624] <= 1'b1;
pika_color[5625] <= 1'b1;
pika_color[5626] <= 1'b1;
pika_color[5627] <= 1'b1;
pika_color[5628] <= 1'b1;
pika_color[5652] <= 1'b1;
pika_color[5670] <= 1'b1;
pika_color[5671] <= 1'b1;
pika_color[5736] <= 1'b1;
pika_color[5737] <= 1'b1;
pika_color[5738] <= 1'b1;
pika_color[5739] <= 1'b1;
pika_color[5740] <= 1'b1;
pika_color[5741] <= 1'b1;
pika_color[5767] <= 1'b1;
pika_color[5768] <= 1'b1;
pika_color[5785] <= 1'b1;
pika_color[5850] <= 1'b1;
pika_color[5851] <= 1'b1;
pika_color[5852] <= 1'b1;
pika_color[5853] <= 1'b1;
pika_color[5854] <= 1'b1;
pika_color[5883] <= 1'b1;
pika_color[5884] <= 1'b1;
pika_color[5899] <= 1'b1;
pika_color[5900] <= 1'b1;
pika_color[5964] <= 1'b1;
pika_color[5965] <= 1'b1;
pika_color[5966] <= 1'b1;
pika_color[5967] <= 1'b1;
pika_color[5999] <= 1'b1;
pika_color[6000] <= 1'b1;
pika_color[6014] <= 1'b1;
pika_color[6076] <= 1'b1;
pika_color[6077] <= 1'b1;
pika_color[6078] <= 1'b1;
pika_color[6079] <= 1'b1;
pika_color[6080] <= 1'b1;
pika_color[6081] <= 1'b1;
pika_color[6115] <= 1'b1;
pika_color[6116] <= 1'b1;
pika_color[6129] <= 1'b1;
pika_color[6176] <= 1'b1;
pika_color[6177] <= 1'b1;
pika_color[6186] <= 1'b1;
pika_color[6187] <= 1'b1;
pika_color[6188] <= 1'b1;
pika_color[6189] <= 1'b1;
pika_color[6190] <= 1'b1;
pika_color[6191] <= 1'b1;
pika_color[6231] <= 1'b1;
pika_color[6232] <= 1'b1;
pika_color[6243] <= 1'b1;
pika_color[6244] <= 1'b1;
pika_color[6292] <= 1'b1;
pika_color[6293] <= 1'b1;
pika_color[6294] <= 1'b1;
pika_color[6295] <= 1'b1;
pika_color[6296] <= 1'b1;
pika_color[6297] <= 1'b1;
pika_color[6298] <= 1'b1;
pika_color[6299] <= 1'b1;
pika_color[6300] <= 1'b1;
pika_color[6301] <= 1'b1;
pika_color[6347] <= 1'b1;
pika_color[6348] <= 1'b1;
pika_color[6358] <= 1'b1;
pika_color[6408] <= 1'b1;
pika_color[6464] <= 1'b1;
pika_color[6472] <= 1'b1;
pika_color[6473] <= 1'b1;
pika_color[6523] <= 1'b1;
pika_color[6580] <= 1'b1;
pika_color[6581] <= 1'b1;
pika_color[6586] <= 1'b1;
pika_color[6587] <= 1'b1;
pika_color[6599] <= 1'b1;
pika_color[6600] <= 1'b1;
pika_color[6638] <= 1'b1;
pika_color[6696] <= 1'b1;
pika_color[6697] <= 1'b1;
pika_color[6701] <= 1'b1;
pika_color[6713] <= 1'b1;
pika_color[6714] <= 1'b1;
pika_color[6715] <= 1'b1;
pika_color[6716] <= 1'b1;
pika_color[6717] <= 1'b1;
pika_color[6753] <= 1'b1;
pika_color[6754] <= 1'b1;
pika_color[6812] <= 1'b1;
pika_color[6816] <= 1'b1;
pika_color[6828] <= 1'b1;
pika_color[6831] <= 1'b1;
pika_color[6832] <= 1'b1;
pika_color[6833] <= 1'b1;
pika_color[6869] <= 1'b1;
pika_color[6927] <= 1'b1;
pika_color[6928] <= 1'b1;
pika_color[6931] <= 1'b1;
pika_color[6942] <= 1'b1;
pika_color[6947] <= 1'b1;
pika_color[6948] <= 1'b1;
pika_color[6949] <= 1'b1;
pika_color[6984] <= 1'b1;
pika_color[7043] <= 1'b1;
pika_color[7046] <= 1'b1;
pika_color[7057] <= 1'b1;
pika_color[7058] <= 1'b1;
pika_color[7061] <= 1'b1;
pika_color[7062] <= 1'b1;
pika_color[7063] <= 1'b1;
pika_color[7064] <= 1'b1;
pika_color[7099] <= 1'b1;
pika_color[7158] <= 1'b1;
pika_color[7161] <= 1'b1;
pika_color[7172] <= 1'b1;
pika_color[7173] <= 1'b1;
pika_color[7174] <= 1'b1;
pika_color[7175] <= 1'b1;
pika_color[7176] <= 1'b1;
pika_color[7177] <= 1'b1;
pika_color[7178] <= 1'b1;
pika_color[7179] <= 1'b1;
pika_color[7200] <= 1'b1;
pika_color[7201] <= 1'b1;
pika_color[7214] <= 1'b1;
pika_color[7273] <= 1'b1;
pika_color[7276] <= 1'b1;
pika_color[7289] <= 1'b1;
pika_color[7290] <= 1'b1;
pika_color[7291] <= 1'b1;
pika_color[7292] <= 1'b1;
pika_color[7293] <= 1'b1;
pika_color[7314] <= 1'b1;
pika_color[7316] <= 1'b1;
pika_color[7317] <= 1'b1;
pika_color[7318] <= 1'b1;
pika_color[7328] <= 1'b1;
pika_color[7389] <= 1'b1;
pika_color[7391] <= 1'b1;
pika_color[7404] <= 1'b1;
pika_color[7405] <= 1'b1;
pika_color[7406] <= 1'b1;
pika_color[7407] <= 1'b1;
pika_color[7428] <= 1'b1;
pika_color[7433] <= 1'b1;
pika_color[7434] <= 1'b1;
pika_color[7443] <= 1'b1;
pika_color[7504] <= 1'b1;
pika_color[7505] <= 1'b1;
pika_color[7543] <= 1'b1;
pika_color[7548] <= 1'b1;
pika_color[7558] <= 1'b1;
pika_color[7618] <= 1'b1;
pika_color[7619] <= 1'b1;
pika_color[7620] <= 1'b1;
pika_color[7658] <= 1'b1;
pika_color[7662] <= 1'b1;
pika_color[7663] <= 1'b1;
pika_color[7664] <= 1'b1;
pika_color[7673] <= 1'b1;
pika_color[7733] <= 1'b1;
pika_color[7735] <= 1'b1;
pika_color[7773] <= 1'b1;
pika_color[7776] <= 1'b1;
pika_color[7777] <= 1'b1;
pika_color[7778] <= 1'b1;
pika_color[7779] <= 1'b1;
pika_color[7788] <= 1'b1;
pika_color[7847] <= 1'b1;
pika_color[7850] <= 1'b1;
pika_color[7890] <= 1'b1;
pika_color[7891] <= 1'b1;
pika_color[7892] <= 1'b1;
pika_color[7893] <= 1'b1;
pika_color[7903] <= 1'b1;
pika_color[7962] <= 1'b1;
pika_color[7966] <= 1'b1;
pika_color[7991] <= 1'b1;
pika_color[7992] <= 1'b1;
pika_color[7993] <= 1'b1;
pika_color[7994] <= 1'b1;
pika_color[8005] <= 1'b1;
pika_color[8006] <= 1'b1;
pika_color[8007] <= 1'b1;
pika_color[8018] <= 1'b1;
pika_color[8076] <= 1'b1;
pika_color[8077] <= 1'b1;
pika_color[8081] <= 1'b1;
pika_color[8106] <= 1'b1;
pika_color[8107] <= 1'b1;
pika_color[8108] <= 1'b1;
pika_color[8109] <= 1'b1;
pika_color[8133] <= 1'b1;
pika_color[8191] <= 1'b1;
pika_color[8196] <= 1'b1;
pika_color[8222] <= 1'b1;
pika_color[8223] <= 1'b1;
pika_color[8248] <= 1'b1;
pika_color[8305] <= 1'b1;
pika_color[8306] <= 1'b1;
pika_color[8310] <= 1'b1;
pika_color[8311] <= 1'b1;
pika_color[8312] <= 1'b1;
pika_color[8362] <= 1'b1;
pika_color[8363] <= 1'b1;
pika_color[8420] <= 1'b1;
pika_color[8425] <= 1'b1;
pika_color[8427] <= 1'b1;
pika_color[8428] <= 1'b1;
pika_color[8477] <= 1'b1;
pika_color[8534] <= 1'b1;
pika_color[8535] <= 1'b1;
pika_color[8539] <= 1'b1;
pika_color[8540] <= 1'b1;
pika_color[8543] <= 1'b1;
pika_color[8592] <= 1'b1;
pika_color[8649] <= 1'b1;
pika_color[8650] <= 1'b1;
pika_color[8654] <= 1'b1;
pika_color[8658] <= 1'b1;
pika_color[8659] <= 1'b1;
pika_color[8681] <= 1'b1;
pika_color[8682] <= 1'b1;
pika_color[8707] <= 1'b1;
pika_color[8765] <= 1'b1;
pika_color[8769] <= 1'b1;
pika_color[8772] <= 1'b1;
pika_color[8773] <= 1'b1;
pika_color[8774] <= 1'b1;
pika_color[8775] <= 1'b1;
pika_color[8776] <= 1'b1;
pika_color[8795] <= 1'b1;
pika_color[8798] <= 1'b1;
pika_color[8821] <= 1'b1;
pika_color[8822] <= 1'b1;
pika_color[8880] <= 1'b1;
pika_color[8881] <= 1'b1;
pika_color[8884] <= 1'b1;
pika_color[8886] <= 1'b1;
pika_color[8887] <= 1'b1;
pika_color[8891] <= 1'b1;
pika_color[8892] <= 1'b1;
pika_color[8893] <= 1'b1;
pika_color[8909] <= 1'b1;
pika_color[8913] <= 1'b1;
pika_color[8936] <= 1'b1;
pika_color[8996] <= 1'b1;
pika_color[8997] <= 1'b1;
pika_color[8998] <= 1'b1;
pika_color[8999] <= 1'b1;
pika_color[9000] <= 1'b1;
pika_color[9008] <= 1'b1;
pika_color[9009] <= 1'b1;
pika_color[9023] <= 1'b1;
pika_color[9028] <= 1'b1;
pika_color[9051] <= 1'b1;
pika_color[9112] <= 1'b1;
pika_color[9113] <= 1'b1;
pika_color[9114] <= 1'b1;
pika_color[9124] <= 1'b1;
pika_color[9138] <= 1'b1;
pika_color[9143] <= 1'b1;
pika_color[9165] <= 1'b1;
pika_color[9166] <= 1'b1;
pika_color[9226] <= 1'b1;
pika_color[9227] <= 1'b1;
pika_color[9228] <= 1'b1;
pika_color[9240] <= 1'b1;
pika_color[9253] <= 1'b1;
pika_color[9258] <= 1'b1;
pika_color[9280] <= 1'b1;
pika_color[9341] <= 1'b1;
pika_color[9355] <= 1'b1;
pika_color[9356] <= 1'b1;
pika_color[9368] <= 1'b1;
pika_color[9373] <= 1'b1;
pika_color[9394] <= 1'b1;
pika_color[9395] <= 1'b1;
pika_color[9455] <= 1'b1;
pika_color[9456] <= 1'b1;
pika_color[9471] <= 1'b1;
pika_color[9472] <= 1'b1;
pika_color[9483] <= 1'b1;
pika_color[9484] <= 1'b1;
pika_color[9485] <= 1'b1;
pika_color[9486] <= 1'b1;
pika_color[9488] <= 1'b1;
pika_color[9509] <= 1'b1;
pika_color[9510] <= 1'b1;
pika_color[9570] <= 1'b1;
pika_color[9587] <= 1'b1;
pika_color[9598] <= 1'b1;
pika_color[9602] <= 1'b1;
pika_color[9603] <= 1'b1;
pika_color[9622] <= 1'b1;
pika_color[9623] <= 1'b1;
pika_color[9625] <= 1'b1;
pika_color[9684] <= 1'b1;
pika_color[9685] <= 1'b1;
pika_color[9703] <= 1'b1;
pika_color[9714] <= 1'b1;
pika_color[9717] <= 1'b1;
pika_color[9735] <= 1'b1;
pika_color[9736] <= 1'b1;
pika_color[9737] <= 1'b1;
pika_color[9741] <= 1'b1;
pika_color[9799] <= 1'b1;
pika_color[9800] <= 1'b1;
pika_color[9818] <= 1'b1;
pika_color[9819] <= 1'b1;
pika_color[9830] <= 1'b1;
pika_color[9831] <= 1'b1;
pika_color[9849] <= 1'b1;
pika_color[9850] <= 1'b1;
pika_color[9856] <= 1'b1;
pika_color[9915] <= 1'b1;
pika_color[9934] <= 1'b1;
pika_color[9963] <= 1'b1;
pika_color[9964] <= 1'b1;
pika_color[9971] <= 1'b1;
pika_color[9972] <= 1'b1;
pika_color[10030] <= 1'b1;
pika_color[10049] <= 1'b1;
pika_color[10050] <= 1'b1;
pika_color[10051] <= 1'b1;
pika_color[10087] <= 1'b1;
pika_color[10145] <= 1'b1;
pika_color[10166] <= 1'b1;
pika_color[10167] <= 1'b1;
pika_color[10202] <= 1'b1;
pika_color[10203] <= 1'b1;
pika_color[10260] <= 1'b1;
pika_color[10282] <= 1'b1;
pika_color[10318] <= 1'b1;
pika_color[10375] <= 1'b1;
pika_color[10398] <= 1'b1;
pika_color[10433] <= 1'b1;
pika_color[10434] <= 1'b1;
pika_color[10489] <= 1'b1;
pika_color[10490] <= 1'b1;
pika_color[10513] <= 1'b1;
pika_color[10549] <= 1'b1;
pika_color[10604] <= 1'b1;
pika_color[10605] <= 1'b1;
pika_color[10606] <= 1'b1;
pika_color[10629] <= 1'b1;
pika_color[10664] <= 1'b1;
pika_color[10665] <= 1'b1;
pika_color[10719] <= 1'b1;
pika_color[10721] <= 1'b1;
pika_color[10722] <= 1'b1;
pika_color[10744] <= 1'b1;
pika_color[10780] <= 1'b1;
pika_color[10834] <= 1'b1;
pika_color[10837] <= 1'b1;
pika_color[10859] <= 1'b1;
pika_color[10860] <= 1'b1;
pika_color[10895] <= 1'b1;
pika_color[10949] <= 1'b1;
pika_color[10952] <= 1'b1;
pika_color[10953] <= 1'b1;
pika_color[10992] <= 1'b1;
pika_color[11010] <= 1'b1;
pika_color[11064] <= 1'b1;
pika_color[11068] <= 1'b1;
pika_color[11069] <= 1'b1;
pika_color[11107] <= 1'b1;
pika_color[11125] <= 1'b1;
pika_color[11126] <= 1'b1;
pika_color[11179] <= 1'b1;
pika_color[11184] <= 1'b1;
pika_color[11222] <= 1'b1;
pika_color[11241] <= 1'b1;
pika_color[11294] <= 1'b1;
pika_color[11338] <= 1'b1;
pika_color[11356] <= 1'b1;
pika_color[11408] <= 1'b1;
pika_color[11409] <= 1'b1;
pika_color[11453] <= 1'b1;
pika_color[11454] <= 1'b1;
pika_color[11471] <= 1'b1;
pika_color[11523] <= 1'b1;
pika_color[11569] <= 1'b1;
pika_color[11586] <= 1'b1;
pika_color[11638] <= 1'b1;
pika_color[11684] <= 1'b1;
pika_color[11685] <= 1'b1;
pika_color[11702] <= 1'b1;
pika_color[11753] <= 1'b1;
pika_color[11800] <= 1'b1;
pika_color[11801] <= 1'b1;
pika_color[11817] <= 1'b1;
pika_color[11868] <= 1'b1;
pika_color[11916] <= 1'b1;
pika_color[11917] <= 1'b1;
pika_color[11932] <= 1'b1;
pika_color[11983] <= 1'b1;
pika_color[12032] <= 1'b1;
pika_color[12047] <= 1'b1;
pika_color[12098] <= 1'b1;
pika_color[12148] <= 1'b1;
pika_color[12162] <= 1'b1;
pika_color[12213] <= 1'b1;
pika_color[12263] <= 1'b1;
pika_color[12264] <= 1'b1;
pika_color[12277] <= 1'b1;
pika_color[12328] <= 1'b1;
pika_color[12379] <= 1'b1;
pika_color[12392] <= 1'b1;
pika_color[12443] <= 1'b1;
pika_color[12494] <= 1'b1;
pika_color[12495] <= 1'b1;
pika_color[12507] <= 1'b1;
pika_color[12558] <= 1'b1;
pika_color[12610] <= 1'b1;
pika_color[12611] <= 1'b1;
pika_color[12621] <= 1'b1;
pika_color[12622] <= 1'b1;
pika_color[12673] <= 1'b1;
pika_color[12727] <= 1'b1;
pika_color[12728] <= 1'b1;
pika_color[12736] <= 1'b1;
pika_color[12788] <= 1'b1;
pika_color[12844] <= 1'b1;
pika_color[12845] <= 1'b1;
pika_color[12851] <= 1'b1;
pika_color[12903] <= 1'b1;
pika_color[12960] <= 1'b1;
pika_color[12961] <= 1'b1;
pika_color[12962] <= 1'b1;
pika_color[12963] <= 1'b1;
pika_color[12964] <= 1'b1;
pika_color[12965] <= 1'b1;
pika_color[13018] <= 1'b1;
pika_color[13077] <= 1'b1;
pika_color[13133] <= 1'b1;
pika_color[13192] <= 1'b1;
pika_color[13248] <= 1'b1;
pika_color[13306] <= 1'b1;
pika_color[13307] <= 1'b1;
pika_color[13363] <= 1'b1;
pika_color[13421] <= 1'b1;
pika_color[13478] <= 1'b1;
pika_color[13536] <= 1'b1;
pika_color[13593] <= 1'b1;
pika_color[13651] <= 1'b1;
pika_color[13708] <= 1'b1;
pika_color[13766] <= 1'b1;
pika_color[13823] <= 1'b1;
pika_color[13824] <= 1'b1;
pika_color[13880] <= 1'b1;
pika_color[13881] <= 1'b1;
pika_color[13939] <= 1'b1;
pika_color[13995] <= 1'b1;
pika_color[14054] <= 1'b1;
pika_color[14055] <= 1'b1;
pika_color[14110] <= 1'b1;
pika_color[14170] <= 1'b1;
pika_color[14171] <= 1'b1;
pika_color[14225] <= 1'b1;
pika_color[14286] <= 1'b1;
pika_color[14339] <= 1'b1;
pika_color[14340] <= 1'b1;
pika_color[14401] <= 1'b1;
pika_color[14454] <= 1'b1;
pika_color[14516] <= 1'b1;
pika_color[14568] <= 1'b1;
pika_color[14569] <= 1'b1;
pika_color[14631] <= 1'b1;
pika_color[14632] <= 1'b1;
pika_color[14682] <= 1'b1;
pika_color[14747] <= 1'b1;
pika_color[14794] <= 1'b1;
pika_color[14795] <= 1'b1;
pika_color[14796] <= 1'b1;
pika_color[14862] <= 1'b1;
pika_color[14863] <= 1'b1;
pika_color[14908] <= 1'b1;
pika_color[14909] <= 1'b1;
pika_color[14978] <= 1'b1;
pika_color[14979] <= 1'b1;
pika_color[15021] <= 1'b1;
pika_color[15022] <= 1'b1;
pika_color[15023] <= 1'b1;
pika_color[15094] <= 1'b1;
pika_color[15095] <= 1'b1;
pika_color[15096] <= 1'b1;
pika_color[15110] <= 1'b1;
pika_color[15111] <= 1'b1;
pika_color[15112] <= 1'b1;
pika_color[15113] <= 1'b1;
pika_color[15114] <= 1'b1;
pika_color[15115] <= 1'b1;
pika_color[15116] <= 1'b1;
pika_color[15117] <= 1'b1;
pika_color[15118] <= 1'b1;
pika_color[15119] <= 1'b1;
pika_color[15120] <= 1'b1;
pika_color[15121] <= 1'b1;
pika_color[15122] <= 1'b1;
pika_color[15123] <= 1'b1;
pika_color[15124] <= 1'b1;
pika_color[15125] <= 1'b1;
pika_color[15126] <= 1'b1;
pika_color[15127] <= 1'b1;
pika_color[15128] <= 1'b1;
pika_color[15129] <= 1'b1;
pika_color[15135] <= 1'b1;
pika_color[15136] <= 1'b1;
pika_color[15137] <= 1'b1;
pika_color[15211] <= 1'b1;
pika_color[15212] <= 1'b1;
pika_color[15224] <= 1'b1;
pika_color[15225] <= 1'b1;
pika_color[15244] <= 1'b1;
pika_color[15245] <= 1'b1;
pika_color[15252] <= 1'b1;
pika_color[15253] <= 1'b1;
pika_color[15327] <= 1'b1;
pika_color[15328] <= 1'b1;
pika_color[15338] <= 1'b1;
pika_color[15339] <= 1'b1;
pika_color[15360] <= 1'b1;
pika_color[15368] <= 1'b1;
pika_color[15369] <= 1'b1;
pika_color[15370] <= 1'b1;
pika_color[15443] <= 1'b1;
pika_color[15453] <= 1'b1;
pika_color[15475] <= 1'b1;
pika_color[15485] <= 1'b1;
pika_color[15559] <= 1'b1;
pika_color[15560] <= 1'b1;
pika_color[15561] <= 1'b1;
pika_color[15562] <= 1'b1;
pika_color[15563] <= 1'b1;
pika_color[15564] <= 1'b1;
pika_color[15565] <= 1'b1;
pika_color[15566] <= 1'b1;
pika_color[15567] <= 1'b1;
pika_color[15568] <= 1'b1;
pika_color[15590] <= 1'b1;
pika_color[15591] <= 1'b1;
pika_color[15599] <= 1'b1;
pika_color[15600] <= 1'b1;
pika_color[15706] <= 1'b1;
pika_color[15707] <= 1'b1;
pika_color[15708] <= 1'b1;
pika_color[15709] <= 1'b1;
pika_color[15710] <= 1'b1;
pika_color[15711] <= 1'b1;
pika_color[15712] <= 1'b1;
pika_color[15713] <= 1'b1;
pika_color[15714] <= 1'b1;

		end
		move10, move11, move12, move13, move14, move15, move16, move17, move18, move19:
		begin
		pika_color[1405] <= 1'b1;
pika_color[1406] <= 1'b1;
pika_color[1519] <= 1'b1;
pika_color[1520] <= 1'b1;
pika_color[1521] <= 1'b1;
pika_color[1522] <= 1'b1;
pika_color[1634] <= 1'b1;
pika_color[1637] <= 1'b1;
pika_color[1638] <= 1'b1;
pika_color[1749] <= 1'b1;
pika_color[1754] <= 1'b1;
pika_color[1864] <= 1'b1;
pika_color[1869] <= 1'b1;
pika_color[1870] <= 1'b1;
pika_color[1978] <= 1'b1;
pika_color[1979] <= 1'b1;
pika_color[1986] <= 1'b1;
pika_color[2093] <= 1'b1;
pika_color[2101] <= 1'b1;
pika_color[2102] <= 1'b1;
pika_color[2196] <= 1'b1;
pika_color[2197] <= 1'b1;
pika_color[2198] <= 1'b1;
pika_color[2199] <= 1'b1;
pika_color[2200] <= 1'b1;
pika_color[2208] <= 1'b1;
pika_color[2217] <= 1'b1;
pika_color[2218] <= 1'b1;
pika_color[2276] <= 1'b1;
pika_color[2277] <= 1'b1;
pika_color[2278] <= 1'b1;
pika_color[2279] <= 1'b1;
pika_color[2310] <= 1'b1;
pika_color[2311] <= 1'b1;
pika_color[2312] <= 1'b1;
pika_color[2313] <= 1'b1;
pika_color[2314] <= 1'b1;
pika_color[2315] <= 1'b1;
pika_color[2316] <= 1'b1;
pika_color[2322] <= 1'b1;
pika_color[2323] <= 1'b1;
pika_color[2333] <= 1'b1;
pika_color[2388] <= 1'b1;
pika_color[2389] <= 1'b1;
pika_color[2390] <= 1'b1;
pika_color[2391] <= 1'b1;
pika_color[2392] <= 1'b1;
pika_color[2393] <= 1'b1;
pika_color[2394] <= 1'b1;
pika_color[2395] <= 1'b1;
pika_color[2396] <= 1'b1;
pika_color[2424] <= 1'b1;
pika_color[2425] <= 1'b1;
pika_color[2426] <= 1'b1;
pika_color[2427] <= 1'b1;
pika_color[2428] <= 1'b1;
pika_color[2429] <= 1'b1;
pika_color[2430] <= 1'b1;
pika_color[2431] <= 1'b1;
pika_color[2432] <= 1'b1;
pika_color[2433] <= 1'b1;
pika_color[2437] <= 1'b1;
pika_color[2448] <= 1'b1;
pika_color[2449] <= 1'b1;
pika_color[2500] <= 1'b1;
pika_color[2501] <= 1'b1;
pika_color[2502] <= 1'b1;
pika_color[2503] <= 1'b1;
pika_color[2506] <= 1'b1;
pika_color[2507] <= 1'b1;
pika_color[2508] <= 1'b1;
pika_color[2509] <= 1'b1;
pika_color[2510] <= 1'b1;
pika_color[2511] <= 1'b1;
pika_color[2512] <= 1'b1;
pika_color[2513] <= 1'b1;
pika_color[2539] <= 1'b1;
pika_color[2540] <= 1'b1;
pika_color[2541] <= 1'b1;
pika_color[2542] <= 1'b1;
pika_color[2543] <= 1'b1;
pika_color[2544] <= 1'b1;
pika_color[2545] <= 1'b1;
pika_color[2548] <= 1'b1;
pika_color[2549] <= 1'b1;
pika_color[2550] <= 1'b1;
pika_color[2551] <= 1'b1;
pika_color[2552] <= 1'b1;
pika_color[2564] <= 1'b1;
pika_color[2565] <= 1'b1;
pika_color[2612] <= 1'b1;
pika_color[2613] <= 1'b1;
pika_color[2614] <= 1'b1;
pika_color[2615] <= 1'b1;
pika_color[2620] <= 1'b1;
pika_color[2621] <= 1'b1;
pika_color[2622] <= 1'b1;
pika_color[2623] <= 1'b1;
pika_color[2624] <= 1'b1;
pika_color[2625] <= 1'b1;
pika_color[2626] <= 1'b1;
pika_color[2627] <= 1'b1;
pika_color[2628] <= 1'b1;
pika_color[2654] <= 1'b1;
pika_color[2655] <= 1'b1;
pika_color[2656] <= 1'b1;
pika_color[2657] <= 1'b1;
pika_color[2658] <= 1'b1;
pika_color[2659] <= 1'b1;
pika_color[2660] <= 1'b1;
pika_color[2666] <= 1'b1;
pika_color[2667] <= 1'b1;
pika_color[2680] <= 1'b1;
pika_color[2726] <= 1'b1;
pika_color[2727] <= 1'b1;
pika_color[2735] <= 1'b1;
pika_color[2736] <= 1'b1;
pika_color[2737] <= 1'b1;
pika_color[2738] <= 1'b1;
pika_color[2739] <= 1'b1;
pika_color[2740] <= 1'b1;
pika_color[2741] <= 1'b1;
pika_color[2742] <= 1'b1;
pika_color[2743] <= 1'b1;
pika_color[2769] <= 1'b1;
pika_color[2770] <= 1'b1;
pika_color[2771] <= 1'b1;
pika_color[2772] <= 1'b1;
pika_color[2773] <= 1'b1;
pika_color[2774] <= 1'b1;
pika_color[2775] <= 1'b1;
pika_color[2782] <= 1'b1;
pika_color[2783] <= 1'b1;
pika_color[2784] <= 1'b1;
pika_color[2785] <= 1'b1;
pika_color[2795] <= 1'b1;
pika_color[2796] <= 1'b1;
pika_color[2839] <= 1'b1;
pika_color[2840] <= 1'b1;
pika_color[2849] <= 1'b1;
pika_color[2850] <= 1'b1;
pika_color[2851] <= 1'b1;
pika_color[2852] <= 1'b1;
pika_color[2853] <= 1'b1;
pika_color[2854] <= 1'b1;
pika_color[2855] <= 1'b1;
pika_color[2856] <= 1'b1;
pika_color[2857] <= 1'b1;
pika_color[2858] <= 1'b1;
pika_color[2884] <= 1'b1;
pika_color[2885] <= 1'b1;
pika_color[2886] <= 1'b1;
pika_color[2887] <= 1'b1;
pika_color[2888] <= 1'b1;
pika_color[2889] <= 1'b1;
pika_color[2890] <= 1'b1;
pika_color[2900] <= 1'b1;
pika_color[2901] <= 1'b1;
pika_color[2902] <= 1'b1;
pika_color[2911] <= 1'b1;
pika_color[2953] <= 1'b1;
pika_color[2954] <= 1'b1;
pika_color[2964] <= 1'b1;
pika_color[2965] <= 1'b1;
pika_color[2966] <= 1'b1;
pika_color[2967] <= 1'b1;
pika_color[2968] <= 1'b1;
pika_color[2969] <= 1'b1;
pika_color[2970] <= 1'b1;
pika_color[2971] <= 1'b1;
pika_color[2972] <= 1'b1;
pika_color[3000] <= 1'b1;
pika_color[3001] <= 1'b1;
pika_color[3002] <= 1'b1;
pika_color[3003] <= 1'b1;
pika_color[3004] <= 1'b1;
pika_color[3005] <= 1'b1;
pika_color[3017] <= 1'b1;
pika_color[3026] <= 1'b1;
pika_color[3027] <= 1'b1;
pika_color[3066] <= 1'b1;
pika_color[3067] <= 1'b1;
pika_color[3068] <= 1'b1;
pika_color[3079] <= 1'b1;
pika_color[3080] <= 1'b1;
pika_color[3081] <= 1'b1;
pika_color[3082] <= 1'b1;
pika_color[3083] <= 1'b1;
pika_color[3084] <= 1'b1;
pika_color[3085] <= 1'b1;
pika_color[3086] <= 1'b1;
pika_color[3087] <= 1'b1;
pika_color[3116] <= 1'b1;
pika_color[3117] <= 1'b1;
pika_color[3118] <= 1'b1;
pika_color[3119] <= 1'b1;
pika_color[3120] <= 1'b1;
pika_color[3133] <= 1'b1;
pika_color[3134] <= 1'b1;
pika_color[3142] <= 1'b1;
pika_color[3180] <= 1'b1;
pika_color[3181] <= 1'b1;
pika_color[3194] <= 1'b1;
pika_color[3195] <= 1'b1;
pika_color[3196] <= 1'b1;
pika_color[3197] <= 1'b1;
pika_color[3198] <= 1'b1;
pika_color[3199] <= 1'b1;
pika_color[3200] <= 1'b1;
pika_color[3201] <= 1'b1;
pika_color[3231] <= 1'b1;
pika_color[3232] <= 1'b1;
pika_color[3233] <= 1'b1;
pika_color[3234] <= 1'b1;
pika_color[3235] <= 1'b1;
pika_color[3249] <= 1'b1;
pika_color[3250] <= 1'b1;
pika_color[3257] <= 1'b1;
pika_color[3258] <= 1'b1;
pika_color[3293] <= 1'b1;
pika_color[3294] <= 1'b1;
pika_color[3308] <= 1'b1;
pika_color[3309] <= 1'b1;
pika_color[3310] <= 1'b1;
pika_color[3311] <= 1'b1;
pika_color[3312] <= 1'b1;
pika_color[3313] <= 1'b1;
pika_color[3314] <= 1'b1;
pika_color[3315] <= 1'b1;
pika_color[3347] <= 1'b1;
pika_color[3348] <= 1'b1;
pika_color[3349] <= 1'b1;
pika_color[3350] <= 1'b1;
pika_color[3365] <= 1'b1;
pika_color[3366] <= 1'b1;
pika_color[3373] <= 1'b1;
pika_color[3407] <= 1'b1;
pika_color[3408] <= 1'b1;
pika_color[3423] <= 1'b1;
pika_color[3424] <= 1'b1;
pika_color[3425] <= 1'b1;
pika_color[3426] <= 1'b1;
pika_color[3427] <= 1'b1;
pika_color[3428] <= 1'b1;
pika_color[3429] <= 1'b1;
pika_color[3462] <= 1'b1;
pika_color[3463] <= 1'b1;
pika_color[3464] <= 1'b1;
pika_color[3465] <= 1'b1;
pika_color[3481] <= 1'b1;
pika_color[3488] <= 1'b1;
pika_color[3489] <= 1'b1;
pika_color[3520] <= 1'b1;
pika_color[3521] <= 1'b1;
pika_color[3522] <= 1'b1;
pika_color[3538] <= 1'b1;
pika_color[3539] <= 1'b1;
pika_color[3540] <= 1'b1;
pika_color[3541] <= 1'b1;
pika_color[3542] <= 1'b1;
pika_color[3543] <= 1'b1;
pika_color[3544] <= 1'b1;
pika_color[3578] <= 1'b1;
pika_color[3579] <= 1'b1;
pika_color[3580] <= 1'b1;
pika_color[3597] <= 1'b1;
pika_color[3598] <= 1'b1;
pika_color[3604] <= 1'b1;
pika_color[3634] <= 1'b1;
pika_color[3635] <= 1'b1;
pika_color[3653] <= 1'b1;
pika_color[3654] <= 1'b1;
pika_color[3655] <= 1'b1;
pika_color[3656] <= 1'b1;
pika_color[3657] <= 1'b1;
pika_color[3658] <= 1'b1;
pika_color[3694] <= 1'b1;
pika_color[3695] <= 1'b1;
pika_color[3713] <= 1'b1;
pika_color[3719] <= 1'b1;
pika_color[3748] <= 1'b1;
pika_color[3749] <= 1'b1;
pika_color[3768] <= 1'b1;
pika_color[3769] <= 1'b1;
pika_color[3770] <= 1'b1;
pika_color[3771] <= 1'b1;
pika_color[3772] <= 1'b1;
pika_color[3810] <= 1'b1;
pika_color[3811] <= 1'b1;
pika_color[3829] <= 1'b1;
pika_color[3834] <= 1'b1;
pika_color[3835] <= 1'b1;
pika_color[3862] <= 1'b1;
pika_color[3863] <= 1'b1;
pika_color[3883] <= 1'b1;
pika_color[3884] <= 1'b1;
pika_color[3885] <= 1'b1;
pika_color[3886] <= 1'b1;
pika_color[3926] <= 1'b1;
pika_color[3944] <= 1'b1;
pika_color[3945] <= 1'b1;
pika_color[3950] <= 1'b1;
pika_color[3959] <= 1'b1;
pika_color[3960] <= 1'b1;
pika_color[3961] <= 1'b1;
pika_color[3962] <= 1'b1;
pika_color[3963] <= 1'b1;
pika_color[3964] <= 1'b1;
pika_color[3965] <= 1'b1;
pika_color[3966] <= 1'b1;
pika_color[3976] <= 1'b1;
pika_color[3977] <= 1'b1;
pika_color[3998] <= 1'b1;
pika_color[3999] <= 1'b1;
pika_color[4041] <= 1'b1;
pika_color[4042] <= 1'b1;
pika_color[4060] <= 1'b1;
pika_color[4061] <= 1'b1;
pika_color[4065] <= 1'b1;
pika_color[4066] <= 1'b1;
pika_color[4069] <= 1'b1;
pika_color[4070] <= 1'b1;
pika_color[4071] <= 1'b1;
pika_color[4072] <= 1'b1;
pika_color[4073] <= 1'b1;
pika_color[4074] <= 1'b1;
pika_color[4081] <= 1'b1;
pika_color[4082] <= 1'b1;
pika_color[4083] <= 1'b1;
pika_color[4084] <= 1'b1;
pika_color[4085] <= 1'b1;
pika_color[4086] <= 1'b1;
pika_color[4090] <= 1'b1;
pika_color[4091] <= 1'b1;
pika_color[4112] <= 1'b1;
pika_color[4113] <= 1'b1;
pika_color[4157] <= 1'b1;
pika_color[4158] <= 1'b1;
pika_color[4176] <= 1'b1;
pika_color[4180] <= 1'b1;
pika_color[4181] <= 1'b1;
pika_color[4182] <= 1'b1;
pika_color[4183] <= 1'b1;
pika_color[4184] <= 1'b1;
pika_color[4201] <= 1'b1;
pika_color[4202] <= 1'b1;
pika_color[4203] <= 1'b1;
pika_color[4204] <= 1'b1;
pika_color[4205] <= 1'b1;
pika_color[4226] <= 1'b1;
pika_color[4227] <= 1'b1;
pika_color[4273] <= 1'b1;
pika_color[4274] <= 1'b1;
pika_color[4291] <= 1'b1;
pika_color[4293] <= 1'b1;
pika_color[4294] <= 1'b1;
pika_color[4295] <= 1'b1;
pika_color[4340] <= 1'b1;
pika_color[4341] <= 1'b1;
pika_color[4389] <= 1'b1;
pika_color[4390] <= 1'b1;
pika_color[4406] <= 1'b1;
pika_color[4407] <= 1'b1;
pika_color[4408] <= 1'b1;
pika_color[4453] <= 1'b1;
pika_color[4454] <= 1'b1;
pika_color[4505] <= 1'b1;
pika_color[4521] <= 1'b1;
pika_color[4522] <= 1'b1;
pika_color[4566] <= 1'b1;
pika_color[4567] <= 1'b1;
pika_color[4620] <= 1'b1;
pika_color[4621] <= 1'b1;
pika_color[4636] <= 1'b1;
pika_color[4637] <= 1'b1;
pika_color[4679] <= 1'b1;
pika_color[4680] <= 1'b1;
pika_color[4681] <= 1'b1;
pika_color[4736] <= 1'b1;
pika_color[4737] <= 1'b1;
pika_color[4791] <= 1'b1;
pika_color[4792] <= 1'b1;
pika_color[4793] <= 1'b1;
pika_color[4794] <= 1'b1;
pika_color[4852] <= 1'b1;
pika_color[4853] <= 1'b1;
pika_color[4904] <= 1'b1;
pika_color[4905] <= 1'b1;
pika_color[4906] <= 1'b1;
pika_color[4968] <= 1'b1;
pika_color[4969] <= 1'b1;
pika_color[5015] <= 1'b1;
pika_color[5016] <= 1'b1;
pika_color[5017] <= 1'b1;
pika_color[5018] <= 1'b1;
pika_color[5084] <= 1'b1;
pika_color[5085] <= 1'b1;
pika_color[5133] <= 1'b1;
pika_color[5134] <= 1'b1;
pika_color[5135] <= 1'b1;
pika_color[5200] <= 1'b1;
pika_color[5201] <= 1'b1;
pika_color[5250] <= 1'b1;
pika_color[5316] <= 1'b1;
pika_color[5317] <= 1'b1;
pika_color[5365] <= 1'b1;
pika_color[5366] <= 1'b1;
pika_color[5432] <= 1'b1;
pika_color[5481] <= 1'b1;
pika_color[5547] <= 1'b1;
pika_color[5548] <= 1'b1;
pika_color[5596] <= 1'b1;
pika_color[5663] <= 1'b1;
pika_color[5664] <= 1'b1;
pika_color[5712] <= 1'b1;
pika_color[5778] <= 1'b1;
pika_color[5827] <= 1'b1;
pika_color[5893] <= 1'b1;
pika_color[5942] <= 1'b1;
pika_color[6008] <= 1'b1;
pika_color[6057] <= 1'b1;
pika_color[6058] <= 1'b1;
pika_color[6122] <= 1'b1;
pika_color[6173] <= 1'b1;
pika_color[6174] <= 1'b1;
pika_color[6237] <= 1'b1;
pika_color[6272] <= 1'b1;
pika_color[6273] <= 1'b1;
pika_color[6274] <= 1'b1;
pika_color[6275] <= 1'b1;
pika_color[6276] <= 1'b1;
pika_color[6288] <= 1'b1;
pika_color[6289] <= 1'b1;
pika_color[6352] <= 1'b1;
pika_color[6386] <= 1'b1;
pika_color[6387] <= 1'b1;
pika_color[6388] <= 1'b1;
pika_color[6389] <= 1'b1;
pika_color[6390] <= 1'b1;
pika_color[6391] <= 1'b1;
pika_color[6392] <= 1'b1;
pika_color[6404] <= 1'b1;
pika_color[6466] <= 1'b1;
pika_color[6467] <= 1'b1;
pika_color[6519] <= 1'b1;
pika_color[6581] <= 1'b1;
pika_color[6592] <= 1'b1;
pika_color[6593] <= 1'b1;
pika_color[6594] <= 1'b1;
pika_color[6595] <= 1'b1;
pika_color[6596] <= 1'b1;
pika_color[6597] <= 1'b1;
pika_color[6598] <= 1'b1;
pika_color[6634] <= 1'b1;
pika_color[6696] <= 1'b1;
pika_color[6706] <= 1'b1;
pika_color[6707] <= 1'b1;
pika_color[6708] <= 1'b1;
pika_color[6709] <= 1'b1;
pika_color[6710] <= 1'b1;
pika_color[6711] <= 1'b1;
pika_color[6712] <= 1'b1;
pika_color[6713] <= 1'b1;
pika_color[6749] <= 1'b1;
pika_color[6811] <= 1'b1;
pika_color[6837] <= 1'b1;
pika_color[6838] <= 1'b1;
pika_color[6839] <= 1'b1;
pika_color[6864] <= 1'b1;
pika_color[6865] <= 1'b1;
pika_color[6866] <= 1'b1;
pika_color[6867] <= 1'b1;
pika_color[6868] <= 1'b1;
pika_color[6869] <= 1'b1;
pika_color[6926] <= 1'b1;
pika_color[6951] <= 1'b1;
pika_color[6952] <= 1'b1;
pika_color[6953] <= 1'b1;
pika_color[6954] <= 1'b1;
pika_color[6977] <= 1'b1;
pika_color[6978] <= 1'b1;
pika_color[6979] <= 1'b1;
pika_color[6984] <= 1'b1;
pika_color[6985] <= 1'b1;
pika_color[6986] <= 1'b1;
pika_color[7041] <= 1'b1;
pika_color[7067] <= 1'b1;
pika_color[7068] <= 1'b1;
pika_color[7092] <= 1'b1;
pika_color[7101] <= 1'b1;
pika_color[7102] <= 1'b1;
pika_color[7156] <= 1'b1;
pika_color[7206] <= 1'b1;
pika_color[7217] <= 1'b1;
pika_color[7271] <= 1'b1;
pika_color[7321] <= 1'b1;
pika_color[7333] <= 1'b1;
pika_color[7386] <= 1'b1;
pika_color[7436] <= 1'b1;
pika_color[7448] <= 1'b1;
pika_color[7449] <= 1'b1;
pika_color[7501] <= 1'b1;
pika_color[7527] <= 1'b1;
pika_color[7528] <= 1'b1;
pika_color[7529] <= 1'b1;
pika_color[7530] <= 1'b1;
pika_color[7531] <= 1'b1;
pika_color[7532] <= 1'b1;
pika_color[7533] <= 1'b1;
pika_color[7551] <= 1'b1;
pika_color[7564] <= 1'b1;
pika_color[7616] <= 1'b1;
pika_color[7639] <= 1'b1;
pika_color[7640] <= 1'b1;
pika_color[7641] <= 1'b1;
pika_color[7642] <= 1'b1;
pika_color[7643] <= 1'b1;
pika_color[7666] <= 1'b1;
pika_color[7679] <= 1'b1;
pika_color[7731] <= 1'b1;
pika_color[7753] <= 1'b1;
pika_color[7754] <= 1'b1;
pika_color[7781] <= 1'b1;
pika_color[7794] <= 1'b1;
pika_color[7846] <= 1'b1;
pika_color[7896] <= 1'b1;
pika_color[7909] <= 1'b1;
pika_color[7962] <= 1'b1;
pika_color[8010] <= 1'b1;
pika_color[8011] <= 1'b1;
pika_color[8024] <= 1'b1;
pika_color[8077] <= 1'b1;
pika_color[8124] <= 1'b1;
pika_color[8125] <= 1'b1;
pika_color[8139] <= 1'b1;
pika_color[8192] <= 1'b1;
pika_color[8238] <= 1'b1;
pika_color[8239] <= 1'b1;
pika_color[8254] <= 1'b1;
pika_color[8307] <= 1'b1;
pika_color[8353] <= 1'b1;
pika_color[8369] <= 1'b1;
pika_color[8423] <= 1'b1;
pika_color[8467] <= 1'b1;
pika_color[8468] <= 1'b1;
pika_color[8484] <= 1'b1;
pika_color[8538] <= 1'b1;
pika_color[8539] <= 1'b1;
pika_color[8582] <= 1'b1;
pika_color[8598] <= 1'b1;
pika_color[8599] <= 1'b1;
pika_color[8654] <= 1'b1;
pika_color[8696] <= 1'b1;
pika_color[8697] <= 1'b1;
pika_color[8712] <= 1'b1;
pika_color[8713] <= 1'b1;
pika_color[8769] <= 1'b1;
pika_color[8770] <= 1'b1;
pika_color[8810] <= 1'b1;
pika_color[8811] <= 1'b1;
pika_color[8827] <= 1'b1;
pika_color[8828] <= 1'b1;
pika_color[8884] <= 1'b1;
pika_color[8885] <= 1'b1;
pika_color[8886] <= 1'b1;
pika_color[8925] <= 1'b1;
pika_color[8942] <= 1'b1;
pika_color[8998] <= 1'b1;
pika_color[8999] <= 1'b1;
pika_color[9001] <= 1'b1;
pika_color[9002] <= 1'b1;
pika_color[9039] <= 1'b1;
pika_color[9040] <= 1'b1;
pika_color[9057] <= 1'b1;
pika_color[9113] <= 1'b1;
pika_color[9118] <= 1'b1;
pika_color[9119] <= 1'b1;
pika_color[9120] <= 1'b1;
pika_color[9153] <= 1'b1;
pika_color[9154] <= 1'b1;
pika_color[9171] <= 1'b1;
pika_color[9228] <= 1'b1;
pika_color[9235] <= 1'b1;
pika_color[9236] <= 1'b1;
pika_color[9237] <= 1'b1;
pika_color[9268] <= 1'b1;
pika_color[9285] <= 1'b1;
pika_color[9286] <= 1'b1;
pika_color[9343] <= 1'b1;
pika_color[9382] <= 1'b1;
pika_color[9383] <= 1'b1;
pika_color[9400] <= 1'b1;
pika_color[9458] <= 1'b1;
pika_color[9496] <= 1'b1;
pika_color[9515] <= 1'b1;
pika_color[9572] <= 1'b1;
pika_color[9573] <= 1'b1;
pika_color[9611] <= 1'b1;
pika_color[9630] <= 1'b1;
pika_color[9687] <= 1'b1;
pika_color[9725] <= 1'b1;
pika_color[9745] <= 1'b1;
pika_color[9802] <= 1'b1;
pika_color[9859] <= 1'b1;
pika_color[9860] <= 1'b1;
pika_color[9917] <= 1'b1;
pika_color[9973] <= 1'b1;
pika_color[9974] <= 1'b1;
pika_color[10032] <= 1'b1;
pika_color[10088] <= 1'b1;
pika_color[10147] <= 1'b1;
pika_color[10202] <= 1'b1;
pika_color[10262] <= 1'b1;
pika_color[10317] <= 1'b1;
pika_color[10377] <= 1'b1;
pika_color[10432] <= 1'b1;
pika_color[10492] <= 1'b1;
pika_color[10547] <= 1'b1;
pika_color[10607] <= 1'b1;
pika_color[10662] <= 1'b1;
pika_color[10663] <= 1'b1;
pika_color[10722] <= 1'b1;
pika_color[10778] <= 1'b1;
pika_color[10837] <= 1'b1;
pika_color[10893] <= 1'b1;
pika_color[10951] <= 1'b1;
pika_color[10952] <= 1'b1;
pika_color[10977] <= 1'b1;
pika_color[11008] <= 1'b1;
pika_color[11066] <= 1'b1;
pika_color[11091] <= 1'b1;
pika_color[11092] <= 1'b1;
pika_color[11123] <= 1'b1;
pika_color[11124] <= 1'b1;
pika_color[11181] <= 1'b1;
pika_color[11206] <= 1'b1;
pika_color[11239] <= 1'b1;
pika_color[11296] <= 1'b1;
pika_color[11320] <= 1'b1;
pika_color[11354] <= 1'b1;
pika_color[11411] <= 1'b1;
pika_color[11434] <= 1'b1;
pika_color[11435] <= 1'b1;
pika_color[11469] <= 1'b1;
pika_color[11526] <= 1'b1;
pika_color[11548] <= 1'b1;
pika_color[11584] <= 1'b1;
pika_color[11641] <= 1'b1;
pika_color[11642] <= 1'b1;
pika_color[11661] <= 1'b1;
pika_color[11662] <= 1'b1;
pika_color[11699] <= 1'b1;
pika_color[11700] <= 1'b1;
pika_color[11756] <= 1'b1;
pika_color[11757] <= 1'b1;
pika_color[11775] <= 1'b1;
pika_color[11776] <= 1'b1;
pika_color[11815] <= 1'b1;
pika_color[11871] <= 1'b1;
pika_color[11872] <= 1'b1;
pika_color[11889] <= 1'b1;
pika_color[11890] <= 1'b1;
pika_color[11930] <= 1'b1;
pika_color[11986] <= 1'b1;
pika_color[11987] <= 1'b1;
pika_color[11988] <= 1'b1;
pika_color[12004] <= 1'b1;
pika_color[12045] <= 1'b1;
pika_color[12100] <= 1'b1;
pika_color[12101] <= 1'b1;
pika_color[12103] <= 1'b1;
pika_color[12119] <= 1'b1;
pika_color[12160] <= 1'b1;
pika_color[12215] <= 1'b1;
pika_color[12218] <= 1'b1;
pika_color[12234] <= 1'b1;
pika_color[12275] <= 1'b1;
pika_color[12330] <= 1'b1;
pika_color[12333] <= 1'b1;
pika_color[12334] <= 1'b1;
pika_color[12349] <= 1'b1;
pika_color[12390] <= 1'b1;
pika_color[12445] <= 1'b1;
pika_color[12449] <= 1'b1;
pika_color[12464] <= 1'b1;
pika_color[12465] <= 1'b1;
pika_color[12505] <= 1'b1;
pika_color[12560] <= 1'b1;
pika_color[12564] <= 1'b1;
pika_color[12565] <= 1'b1;
pika_color[12580] <= 1'b1;
pika_color[12620] <= 1'b1;
pika_color[12675] <= 1'b1;
pika_color[12680] <= 1'b1;
pika_color[12695] <= 1'b1;
pika_color[12735] <= 1'b1;
pika_color[12790] <= 1'b1;
pika_color[12795] <= 1'b1;
pika_color[12809] <= 1'b1;
pika_color[12810] <= 1'b1;
pika_color[12850] <= 1'b1;
pika_color[12905] <= 1'b1;
pika_color[12910] <= 1'b1;
pika_color[12911] <= 1'b1;
pika_color[12924] <= 1'b1;
pika_color[12964] <= 1'b1;
pika_color[12965] <= 1'b1;
pika_color[13020] <= 1'b1;
pika_color[13026] <= 1'b1;
pika_color[13038] <= 1'b1;
pika_color[13079] <= 1'b1;
pika_color[13135] <= 1'b1;
pika_color[13136] <= 1'b1;
pika_color[13142] <= 1'b1;
pika_color[13152] <= 1'b1;
pika_color[13153] <= 1'b1;
pika_color[13194] <= 1'b1;
pika_color[13251] <= 1'b1;
pika_color[13258] <= 1'b1;
pika_color[13259] <= 1'b1;
pika_color[13266] <= 1'b1;
pika_color[13267] <= 1'b1;
pika_color[13309] <= 1'b1;
pika_color[13366] <= 1'b1;
pika_color[13374] <= 1'b1;
pika_color[13375] <= 1'b1;
pika_color[13376] <= 1'b1;
pika_color[13377] <= 1'b1;
pika_color[13378] <= 1'b1;
pika_color[13379] <= 1'b1;
pika_color[13380] <= 1'b1;
pika_color[13381] <= 1'b1;
pika_color[13424] <= 1'b1;
pika_color[13481] <= 1'b1;
pika_color[13539] <= 1'b1;
pika_color[13596] <= 1'b1;
pika_color[13597] <= 1'b1;
pika_color[13654] <= 1'b1;
pika_color[13712] <= 1'b1;
pika_color[13768] <= 1'b1;
pika_color[13769] <= 1'b1;
pika_color[13827] <= 1'b1;
pika_color[13883] <= 1'b1;
pika_color[13942] <= 1'b1;
pika_color[13998] <= 1'b1;
pika_color[14057] <= 1'b1;
pika_color[14058] <= 1'b1;
pika_color[14112] <= 1'b1;
pika_color[14173] <= 1'b1;
pika_color[14226] <= 1'b1;
pika_color[14227] <= 1'b1;
pika_color[14288] <= 1'b1;
pika_color[14289] <= 1'b1;
pika_color[14340] <= 1'b1;
pika_color[14341] <= 1'b1;
pika_color[14404] <= 1'b1;
pika_color[14454] <= 1'b1;
pika_color[14455] <= 1'b1;
pika_color[14519] <= 1'b1;
pika_color[14520] <= 1'b1;
pika_color[14569] <= 1'b1;
pika_color[14635] <= 1'b1;
pika_color[14683] <= 1'b1;
pika_color[14684] <= 1'b1;
pika_color[14750] <= 1'b1;
pika_color[14751] <= 1'b1;
pika_color[14797] <= 1'b1;
pika_color[14798] <= 1'b1;
pika_color[14866] <= 1'b1;
pika_color[14867] <= 1'b1;
pika_color[14911] <= 1'b1;
pika_color[14912] <= 1'b1;
pika_color[14982] <= 1'b1;
pika_color[14983] <= 1'b1;
pika_color[15002] <= 1'b1;
pika_color[15003] <= 1'b1;
pika_color[15004] <= 1'b1;
pika_color[15005] <= 1'b1;
pika_color[15006] <= 1'b1;
pika_color[15007] <= 1'b1;
pika_color[15008] <= 1'b1;
pika_color[15009] <= 1'b1;
pika_color[15025] <= 1'b1;
pika_color[15026] <= 1'b1;
pika_color[15098] <= 1'b1;
pika_color[15099] <= 1'b1;
pika_color[15100] <= 1'b1;
pika_color[15115] <= 1'b1;
pika_color[15116] <= 1'b1;
pika_color[15117] <= 1'b1;
pika_color[15124] <= 1'b1;
pika_color[15125] <= 1'b1;
pika_color[15138] <= 1'b1;
pika_color[15139] <= 1'b1;
pika_color[15140] <= 1'b1;
pika_color[15215] <= 1'b1;
pika_color[15216] <= 1'b1;
pika_color[15217] <= 1'b1;
pika_color[15218] <= 1'b1;
pika_color[15229] <= 1'b1;
pika_color[15230] <= 1'b1;
pika_color[15240] <= 1'b1;
pika_color[15241] <= 1'b1;
pika_color[15242] <= 1'b1;
pika_color[15252] <= 1'b1;
pika_color[15253] <= 1'b1;
pika_color[15333] <= 1'b1;
pika_color[15334] <= 1'b1;
pika_color[15335] <= 1'b1;
pika_color[15336] <= 1'b1;
pika_color[15337] <= 1'b1;
pika_color[15338] <= 1'b1;
pika_color[15339] <= 1'b1;
pika_color[15345] <= 1'b1;
pika_color[15346] <= 1'b1;
pika_color[15357] <= 1'b1;
pika_color[15358] <= 1'b1;
pika_color[15359] <= 1'b1;
pika_color[15360] <= 1'b1;
pika_color[15361] <= 1'b1;
pika_color[15362] <= 1'b1;
pika_color[15363] <= 1'b1;
pika_color[15364] <= 1'b1;
pika_color[15365] <= 1'b1;
pika_color[15366] <= 1'b1;
pika_color[15452] <= 1'b1;
pika_color[15453] <= 1'b1;
pika_color[15461] <= 1'b1;
pika_color[15462] <= 1'b1;
pika_color[15567] <= 1'b1;
pika_color[15577] <= 1'b1;
pika_color[15682] <= 1'b1;
pika_color[15692] <= 1'b1;
pika_color[15797] <= 1'b1;
pika_color[15799] <= 1'b1;
pika_color[15800] <= 1'b1;
pika_color[15801] <= 1'b1;
pika_color[15802] <= 1'b1;
pika_color[15803] <= 1'b1;
pika_color[15804] <= 1'b1;
pika_color[15805] <= 1'b1;
pika_color[15806] <= 1'b1;
pika_color[15807] <= 1'b1;
pika_color[15912] <= 1'b1;
pika_color[15913] <= 1'b1;
pika_color[15914] <= 1'b1;

		end
		move20, move21, move22, move23, move24, move25, move26, move27, move28, move29:
		begin
		
pika_color[1852] <= 1'b1;
pika_color[1853] <= 1'b1;
pika_color[1854] <= 1'b1;
pika_color[1966] <= 1'b1;
pika_color[1967] <= 1'b1;
pika_color[1968] <= 1'b1;
pika_color[1969] <= 1'b1;
pika_color[1970] <= 1'b1;
pika_color[2081] <= 1'b1;
pika_color[2082] <= 1'b1;
pika_color[2083] <= 1'b1;
pika_color[2084] <= 1'b1;
pika_color[2085] <= 1'b1;
pika_color[2086] <= 1'b1;
pika_color[2150] <= 1'b1;
pika_color[2151] <= 1'b1;
pika_color[2152] <= 1'b1;
pika_color[2153] <= 1'b1;
pika_color[2154] <= 1'b1;
pika_color[2155] <= 1'b1;
pika_color[2196] <= 1'b1;
pika_color[2197] <= 1'b1;
pika_color[2198] <= 1'b1;
pika_color[2199] <= 1'b1;
pika_color[2200] <= 1'b1;
pika_color[2201] <= 1'b1;
pika_color[2202] <= 1'b1;
pika_color[2203] <= 1'b1;
pika_color[2263] <= 1'b1;
pika_color[2264] <= 1'b1;
pika_color[2265] <= 1'b1;
pika_color[2266] <= 1'b1;
pika_color[2267] <= 1'b1;
pika_color[2268] <= 1'b1;
pika_color[2269] <= 1'b1;
pika_color[2270] <= 1'b1;
pika_color[2310] <= 1'b1;
pika_color[2311] <= 1'b1;
pika_color[2312] <= 1'b1;
pika_color[2313] <= 1'b1;
pika_color[2314] <= 1'b1;
pika_color[2315] <= 1'b1;
pika_color[2316] <= 1'b1;
pika_color[2317] <= 1'b1;
pika_color[2318] <= 1'b1;
pika_color[2319] <= 1'b1;
pika_color[2376] <= 1'b1;
pika_color[2377] <= 1'b1;
pika_color[2378] <= 1'b1;
pika_color[2379] <= 1'b1;
pika_color[2380] <= 1'b1;
pika_color[2381] <= 1'b1;
pika_color[2382] <= 1'b1;
pika_color[2383] <= 1'b1;
pika_color[2384] <= 1'b1;
pika_color[2385] <= 1'b1;
pika_color[2425] <= 1'b1;
pika_color[2426] <= 1'b1;
pika_color[2427] <= 1'b1;
pika_color[2428] <= 1'b1;
pika_color[2429] <= 1'b1;
pika_color[2430] <= 1'b1;
pika_color[2431] <= 1'b1;
pika_color[2432] <= 1'b1;
pika_color[2433] <= 1'b1;
pika_color[2434] <= 1'b1;
pika_color[2490] <= 1'b1;
pika_color[2491] <= 1'b1;
pika_color[2494] <= 1'b1;
pika_color[2495] <= 1'b1;
pika_color[2496] <= 1'b1;
pika_color[2497] <= 1'b1;
pika_color[2498] <= 1'b1;
pika_color[2499] <= 1'b1;
pika_color[2500] <= 1'b1;
pika_color[2540] <= 1'b1;
pika_color[2541] <= 1'b1;
pika_color[2542] <= 1'b1;
pika_color[2543] <= 1'b1;
pika_color[2544] <= 1'b1;
pika_color[2545] <= 1'b1;
pika_color[2546] <= 1'b1;
pika_color[2547] <= 1'b1;
pika_color[2549] <= 1'b1;
pika_color[2550] <= 1'b1;
pika_color[2604] <= 1'b1;
pika_color[2605] <= 1'b1;
pika_color[2609] <= 1'b1;
pika_color[2610] <= 1'b1;
pika_color[2611] <= 1'b1;
pika_color[2612] <= 1'b1;
pika_color[2613] <= 1'b1;
pika_color[2614] <= 1'b1;
pika_color[2615] <= 1'b1;
pika_color[2655] <= 1'b1;
pika_color[2656] <= 1'b1;
pika_color[2657] <= 1'b1;
pika_color[2658] <= 1'b1;
pika_color[2659] <= 1'b1;
pika_color[2660] <= 1'b1;
pika_color[2661] <= 1'b1;
pika_color[2662] <= 1'b1;
pika_color[2665] <= 1'b1;
pika_color[2666] <= 1'b1;
pika_color[2718] <= 1'b1;
pika_color[2719] <= 1'b1;
pika_color[2724] <= 1'b1;
pika_color[2725] <= 1'b1;
pika_color[2726] <= 1'b1;
pika_color[2727] <= 1'b1;
pika_color[2728] <= 1'b1;
pika_color[2729] <= 1'b1;
pika_color[2770] <= 1'b1;
pika_color[2771] <= 1'b1;
pika_color[2772] <= 1'b1;
pika_color[2773] <= 1'b1;
pika_color[2774] <= 1'b1;
pika_color[2775] <= 1'b1;
pika_color[2776] <= 1'b1;
pika_color[2781] <= 1'b1;
pika_color[2782] <= 1'b1;
pika_color[2832] <= 1'b1;
pika_color[2833] <= 1'b1;
pika_color[2839] <= 1'b1;
pika_color[2840] <= 1'b1;
pika_color[2841] <= 1'b1;
pika_color[2842] <= 1'b1;
pika_color[2843] <= 1'b1;
pika_color[2844] <= 1'b1;
pika_color[2885] <= 1'b1;
pika_color[2886] <= 1'b1;
pika_color[2887] <= 1'b1;
pika_color[2888] <= 1'b1;
pika_color[2889] <= 1'b1;
pika_color[2890] <= 1'b1;
pika_color[2891] <= 1'b1;
pika_color[2897] <= 1'b1;
pika_color[2946] <= 1'b1;
pika_color[2947] <= 1'b1;
pika_color[2954] <= 1'b1;
pika_color[2955] <= 1'b1;
pika_color[2956] <= 1'b1;
pika_color[2957] <= 1'b1;
pika_color[2958] <= 1'b1;
pika_color[2959] <= 1'b1;
pika_color[3001] <= 1'b1;
pika_color[3002] <= 1'b1;
pika_color[3003] <= 1'b1;
pika_color[3004] <= 1'b1;
pika_color[3005] <= 1'b1;
pika_color[3012] <= 1'b1;
pika_color[3013] <= 1'b1;
pika_color[3060] <= 1'b1;
pika_color[3061] <= 1'b1;
pika_color[3069] <= 1'b1;
pika_color[3070] <= 1'b1;
pika_color[3071] <= 1'b1;
pika_color[3072] <= 1'b1;
pika_color[3073] <= 1'b1;
pika_color[3074] <= 1'b1;
pika_color[3116] <= 1'b1;
pika_color[3117] <= 1'b1;
pika_color[3118] <= 1'b1;
pika_color[3119] <= 1'b1;
pika_color[3120] <= 1'b1;
pika_color[3128] <= 1'b1;
pika_color[3129] <= 1'b1;
pika_color[3174] <= 1'b1;
pika_color[3175] <= 1'b1;
pika_color[3184] <= 1'b1;
pika_color[3185] <= 1'b1;
pika_color[3186] <= 1'b1;
pika_color[3187] <= 1'b1;
pika_color[3188] <= 1'b1;
pika_color[3231] <= 1'b1;
pika_color[3232] <= 1'b1;
pika_color[3233] <= 1'b1;
pika_color[3234] <= 1'b1;
pika_color[3244] <= 1'b1;
pika_color[3288] <= 1'b1;
pika_color[3289] <= 1'b1;
pika_color[3299] <= 1'b1;
pika_color[3300] <= 1'b1;
pika_color[3301] <= 1'b1;
pika_color[3302] <= 1'b1;
pika_color[3303] <= 1'b1;
pika_color[3346] <= 1'b1;
pika_color[3347] <= 1'b1;
pika_color[3348] <= 1'b1;
pika_color[3349] <= 1'b1;
pika_color[3359] <= 1'b1;
pika_color[3360] <= 1'b1;
pika_color[3402] <= 1'b1;
pika_color[3403] <= 1'b1;
pika_color[3415] <= 1'b1;
pika_color[3416] <= 1'b1;
pika_color[3417] <= 1'b1;
pika_color[3462] <= 1'b1;
pika_color[3463] <= 1'b1;
pika_color[3475] <= 1'b1;
pika_color[3476] <= 1'b1;
pika_color[3516] <= 1'b1;
pika_color[3517] <= 1'b1;
pika_color[3530] <= 1'b1;
pika_color[3531] <= 1'b1;
pika_color[3532] <= 1'b1;
pika_color[3577] <= 1'b1;
pika_color[3578] <= 1'b1;
pika_color[3591] <= 1'b1;
pika_color[3630] <= 1'b1;
pika_color[3631] <= 1'b1;
pika_color[3645] <= 1'b1;
pika_color[3646] <= 1'b1;
pika_color[3647] <= 1'b1;
pika_color[3692] <= 1'b1;
pika_color[3693] <= 1'b1;
pika_color[3706] <= 1'b1;
pika_color[3707] <= 1'b1;
pika_color[3745] <= 1'b1;
pika_color[3760] <= 1'b1;
pika_color[3761] <= 1'b1;
pika_color[3807] <= 1'b1;
pika_color[3808] <= 1'b1;
pika_color[3822] <= 1'b1;
pika_color[3859] <= 1'b1;
pika_color[3875] <= 1'b1;
pika_color[3876] <= 1'b1;
pika_color[3923] <= 1'b1;
pika_color[3924] <= 1'b1;
pika_color[3937] <= 1'b1;
pika_color[3974] <= 1'b1;
pika_color[3990] <= 1'b1;
pika_color[3991] <= 1'b1;
pika_color[4038] <= 1'b1;
pika_color[4039] <= 1'b1;
pika_color[4052] <= 1'b1;
pika_color[4053] <= 1'b1;
pika_color[4088] <= 1'b1;
pika_color[4089] <= 1'b1;
pika_color[4105] <= 1'b1;
pika_color[4154] <= 1'b1;
pika_color[4168] <= 1'b1;
pika_color[4169] <= 1'b1;
pika_color[4203] <= 1'b1;
pika_color[4219] <= 1'b1;
pika_color[4220] <= 1'b1;
pika_color[4269] <= 1'b1;
pika_color[4270] <= 1'b1;
pika_color[4284] <= 1'b1;
pika_color[4317] <= 1'b1;
pika_color[4318] <= 1'b1;
pika_color[4334] <= 1'b1;
pika_color[4385] <= 1'b1;
pika_color[4399] <= 1'b1;
pika_color[4432] <= 1'b1;
pika_color[4448] <= 1'b1;
pika_color[4449] <= 1'b1;
pika_color[4500] <= 1'b1;
pika_color[4514] <= 1'b1;
pika_color[4515] <= 1'b1;
pika_color[4546] <= 1'b1;
pika_color[4547] <= 1'b1;
pika_color[4563] <= 1'b1;
pika_color[4615] <= 1'b1;
pika_color[4616] <= 1'b1;
pika_color[4630] <= 1'b1;
pika_color[4661] <= 1'b1;
pika_color[4677] <= 1'b1;
pika_color[4678] <= 1'b1;
pika_color[4725] <= 1'b1;
pika_color[4726] <= 1'b1;
pika_color[4727] <= 1'b1;
pika_color[4731] <= 1'b1;
pika_color[4745] <= 1'b1;
pika_color[4746] <= 1'b1;
pika_color[4776] <= 1'b1;
pika_color[4791] <= 1'b1;
pika_color[4839] <= 1'b1;
pika_color[4840] <= 1'b1;
pika_color[4842] <= 1'b1;
pika_color[4843] <= 1'b1;
pika_color[4846] <= 1'b1;
pika_color[4861] <= 1'b1;
pika_color[4873] <= 1'b1;
pika_color[4874] <= 1'b1;
pika_color[4875] <= 1'b1;
pika_color[4876] <= 1'b1;
pika_color[4877] <= 1'b1;
pika_color[4878] <= 1'b1;
pika_color[4879] <= 1'b1;
pika_color[4890] <= 1'b1;
pika_color[4905] <= 1'b1;
pika_color[4906] <= 1'b1;
pika_color[4953] <= 1'b1;
pika_color[4954] <= 1'b1;
pika_color[4959] <= 1'b1;
pika_color[4961] <= 1'b1;
pika_color[4976] <= 1'b1;
pika_color[4981] <= 1'b1;
pika_color[4982] <= 1'b1;
pika_color[4983] <= 1'b1;
pika_color[4984] <= 1'b1;
pika_color[4985] <= 1'b1;
pika_color[4986] <= 1'b1;
pika_color[4987] <= 1'b1;
pika_color[4995] <= 1'b1;
pika_color[4996] <= 1'b1;
pika_color[4997] <= 1'b1;
pika_color[4998] <= 1'b1;
pika_color[5004] <= 1'b1;
pika_color[5005] <= 1'b1;
pika_color[5019] <= 1'b1;
pika_color[5020] <= 1'b1;
pika_color[5068] <= 1'b1;
pika_color[5074] <= 1'b1;
pika_color[5075] <= 1'b1;
pika_color[5076] <= 1'b1;
pika_color[5077] <= 1'b1;
pika_color[5091] <= 1'b1;
pika_color[5092] <= 1'b1;
pika_color[5094] <= 1'b1;
pika_color[5095] <= 1'b1;
pika_color[5096] <= 1'b1;
pika_color[5113] <= 1'b1;
pika_color[5114] <= 1'b1;
pika_color[5115] <= 1'b1;
pika_color[5116] <= 1'b1;
pika_color[5119] <= 1'b1;
pika_color[5133] <= 1'b1;
pika_color[5134] <= 1'b1;
pika_color[5183] <= 1'b1;
pika_color[5190] <= 1'b1;
pika_color[5191] <= 1'b1;
pika_color[5192] <= 1'b1;
pika_color[5206] <= 1'b1;
pika_color[5207] <= 1'b1;
pika_color[5208] <= 1'b1;
pika_color[5209] <= 1'b1;
pika_color[5231] <= 1'b1;
pika_color[5232] <= 1'b1;
pika_color[5233] <= 1'b1;
pika_color[5234] <= 1'b1;
pika_color[5247] <= 1'b1;
pika_color[5248] <= 1'b1;
pika_color[5298] <= 1'b1;
pika_color[5306] <= 1'b1;
pika_color[5307] <= 1'b1;
pika_color[5308] <= 1'b1;
pika_color[5322] <= 1'b1;
pika_color[5361] <= 1'b1;
pika_color[5362] <= 1'b1;
pika_color[5413] <= 1'b1;
pika_color[5422] <= 1'b1;
pika_color[5423] <= 1'b1;
pika_color[5475] <= 1'b1;
pika_color[5476] <= 1'b1;
pika_color[5528] <= 1'b1;
pika_color[5538] <= 1'b1;
pika_color[5539] <= 1'b1;
pika_color[5589] <= 1'b1;
pika_color[5590] <= 1'b1;
pika_color[5643] <= 1'b1;
pika_color[5653] <= 1'b1;
pika_color[5654] <= 1'b1;
pika_color[5655] <= 1'b1;
pika_color[5703] <= 1'b1;
pika_color[5704] <= 1'b1;
pika_color[5758] <= 1'b1;
pika_color[5769] <= 1'b1;
pika_color[5770] <= 1'b1;
pika_color[5817] <= 1'b1;
pika_color[5818] <= 1'b1;
pika_color[5873] <= 1'b1;
pika_color[5884] <= 1'b1;
pika_color[5885] <= 1'b1;
pika_color[5931] <= 1'b1;
pika_color[5932] <= 1'b1;
pika_color[5988] <= 1'b1;
pika_color[6000] <= 1'b1;
pika_color[6001] <= 1'b1;
pika_color[6046] <= 1'b1;
pika_color[6047] <= 1'b1;
pika_color[6103] <= 1'b1;
pika_color[6115] <= 1'b1;
pika_color[6116] <= 1'b1;
pika_color[6162] <= 1'b1;
pika_color[6163] <= 1'b1;
pika_color[6218] <= 1'b1;
pika_color[6231] <= 1'b1;
pika_color[6278] <= 1'b1;
pika_color[6279] <= 1'b1;
pika_color[6333] <= 1'b1;
pika_color[6346] <= 1'b1;
pika_color[6347] <= 1'b1;
pika_color[6394] <= 1'b1;
pika_color[6448] <= 1'b1;
pika_color[6449] <= 1'b1;
pika_color[6462] <= 1'b1;
pika_color[6509] <= 1'b1;
pika_color[6564] <= 1'b1;
pika_color[6578] <= 1'b1;
pika_color[6625] <= 1'b1;
pika_color[6679] <= 1'b1;
pika_color[6693] <= 1'b1;
pika_color[6694] <= 1'b1;
pika_color[6740] <= 1'b1;
pika_color[6794] <= 1'b1;
pika_color[6808] <= 1'b1;
pika_color[6855] <= 1'b1;
pika_color[6909] <= 1'b1;
pika_color[6922] <= 1'b1;
pika_color[6923] <= 1'b1;
pika_color[6970] <= 1'b1;
pika_color[6971] <= 1'b1;
pika_color[7024] <= 1'b1;
pika_color[7037] <= 1'b1;
pika_color[7086] <= 1'b1;
pika_color[7139] <= 1'b1;
pika_color[7152] <= 1'b1;
pika_color[7201] <= 1'b1;
pika_color[7254] <= 1'b1;
pika_color[7267] <= 1'b1;
pika_color[7316] <= 1'b1;
pika_color[7369] <= 1'b1;
pika_color[7370] <= 1'b1;
pika_color[7382] <= 1'b1;
pika_color[7431] <= 1'b1;
pika_color[7485] <= 1'b1;
pika_color[7496] <= 1'b1;
pika_color[7546] <= 1'b1;
pika_color[7547] <= 1'b1;
pika_color[7600] <= 1'b1;
pika_color[7611] <= 1'b1;
pika_color[7646] <= 1'b1;
pika_color[7647] <= 1'b1;
pika_color[7648] <= 1'b1;
pika_color[7649] <= 1'b1;
pika_color[7650] <= 1'b1;
pika_color[7662] <= 1'b1;
pika_color[7715] <= 1'b1;
pika_color[7726] <= 1'b1;
pika_color[7760] <= 1'b1;
pika_color[7761] <= 1'b1;
pika_color[7762] <= 1'b1;
pika_color[7763] <= 1'b1;
pika_color[7764] <= 1'b1;
pika_color[7777] <= 1'b1;
pika_color[7778] <= 1'b1;
pika_color[7830] <= 1'b1;
pika_color[7841] <= 1'b1;
pika_color[7890] <= 1'b1;
pika_color[7891] <= 1'b1;
pika_color[7892] <= 1'b1;
pika_color[7893] <= 1'b1;
pika_color[7945] <= 1'b1;
pika_color[7946] <= 1'b1;
pika_color[7956] <= 1'b1;
pika_color[7966] <= 1'b1;
pika_color[7967] <= 1'b1;
pika_color[7968] <= 1'b1;
pika_color[7969] <= 1'b1;
pika_color[7970] <= 1'b1;
pika_color[7971] <= 1'b1;
pika_color[7972] <= 1'b1;
pika_color[8003] <= 1'b1;
pika_color[8004] <= 1'b1;
pika_color[8005] <= 1'b1;
pika_color[8008] <= 1'b1;
pika_color[8009] <= 1'b1;
pika_color[8010] <= 1'b1;
pika_color[8011] <= 1'b1;
pika_color[8061] <= 1'b1;
pika_color[8071] <= 1'b1;
pika_color[8082] <= 1'b1;
pika_color[8083] <= 1'b1;
pika_color[8084] <= 1'b1;
pika_color[8085] <= 1'b1;
pika_color[8086] <= 1'b1;
pika_color[8087] <= 1'b1;
pika_color[8116] <= 1'b1;
pika_color[8117] <= 1'b1;
pika_color[8118] <= 1'b1;
pika_color[8126] <= 1'b1;
pika_color[8127] <= 1'b1;
pika_color[8176] <= 1'b1;
pika_color[8186] <= 1'b1;
pika_color[8230] <= 1'b1;
pika_color[8231] <= 1'b1;
pika_color[8242] <= 1'b1;
pika_color[8243] <= 1'b1;
pika_color[8291] <= 1'b1;
pika_color[8292] <= 1'b1;
pika_color[8301] <= 1'b1;
pika_color[8345] <= 1'b1;
pika_color[8358] <= 1'b1;
pika_color[8407] <= 1'b1;
pika_color[8416] <= 1'b1;
pika_color[8440] <= 1'b1;
pika_color[8441] <= 1'b1;
pika_color[8442] <= 1'b1;
pika_color[8443] <= 1'b1;
pika_color[8444] <= 1'b1;
pika_color[8460] <= 1'b1;
pika_color[8473] <= 1'b1;
pika_color[8522] <= 1'b1;
pika_color[8531] <= 1'b1;
pika_color[8556] <= 1'b1;
pika_color[8557] <= 1'b1;
pika_color[8558] <= 1'b1;
pika_color[8575] <= 1'b1;
pika_color[8588] <= 1'b1;
pika_color[8637] <= 1'b1;
pika_color[8638] <= 1'b1;
pika_color[8646] <= 1'b1;
pika_color[8690] <= 1'b1;
pika_color[8703] <= 1'b1;
pika_color[8753] <= 1'b1;
pika_color[8754] <= 1'b1;
pika_color[8755] <= 1'b1;
pika_color[8761] <= 1'b1;
pika_color[8805] <= 1'b1;
pika_color[8818] <= 1'b1;
pika_color[8870] <= 1'b1;
pika_color[8871] <= 1'b1;
pika_color[8872] <= 1'b1;
pika_color[8873] <= 1'b1;
pika_color[8874] <= 1'b1;
pika_color[8875] <= 1'b1;
pika_color[8876] <= 1'b1;
pika_color[8920] <= 1'b1;
pika_color[8933] <= 1'b1;
pika_color[8990] <= 1'b1;
pika_color[8991] <= 1'b1;
pika_color[9035] <= 1'b1;
pika_color[9048] <= 1'b1;
pika_color[9106] <= 1'b1;
pika_color[9131] <= 1'b1;
pika_color[9132] <= 1'b1;
pika_color[9133] <= 1'b1;
pika_color[9134] <= 1'b1;
pika_color[9150] <= 1'b1;
pika_color[9163] <= 1'b1;
pika_color[9221] <= 1'b1;
pika_color[9244] <= 1'b1;
pika_color[9245] <= 1'b1;
pika_color[9250] <= 1'b1;
pika_color[9251] <= 1'b1;
pika_color[9252] <= 1'b1;
pika_color[9265] <= 1'b1;
pika_color[9278] <= 1'b1;
pika_color[9336] <= 1'b1;
pika_color[9337] <= 1'b1;
pika_color[9357] <= 1'b1;
pika_color[9358] <= 1'b1;
pika_color[9359] <= 1'b1;
pika_color[9368] <= 1'b1;
pika_color[9380] <= 1'b1;
pika_color[9393] <= 1'b1;
pika_color[9452] <= 1'b1;
pika_color[9472] <= 1'b1;
pika_color[9483] <= 1'b1;
pika_color[9495] <= 1'b1;
pika_color[9508] <= 1'b1;
pika_color[9568] <= 1'b1;
pika_color[9588] <= 1'b1;
pika_color[9597] <= 1'b1;
pika_color[9598] <= 1'b1;
pika_color[9610] <= 1'b1;
pika_color[9623] <= 1'b1;
pika_color[9683] <= 1'b1;
pika_color[9684] <= 1'b1;
pika_color[9703] <= 1'b1;
pika_color[9706] <= 1'b1;
pika_color[9707] <= 1'b1;
pika_color[9708] <= 1'b1;
pika_color[9709] <= 1'b1;
pika_color[9710] <= 1'b1;
pika_color[9712] <= 1'b1;
pika_color[9725] <= 1'b1;
pika_color[9738] <= 1'b1;
pika_color[9797] <= 1'b1;
pika_color[9798] <= 1'b1;
pika_color[9799] <= 1'b1;
pika_color[9818] <= 1'b1;
pika_color[9819] <= 1'b1;
pika_color[9820] <= 1'b1;
pika_color[9821] <= 1'b1;
pika_color[9825] <= 1'b1;
pika_color[9826] <= 1'b1;
pika_color[9827] <= 1'b1;
pika_color[9840] <= 1'b1;
pika_color[9853] <= 1'b1;
pika_color[9911] <= 1'b1;
pika_color[9912] <= 1'b1;
pika_color[9914] <= 1'b1;
pika_color[9915] <= 1'b1;
pika_color[9934] <= 1'b1;
pika_color[9941] <= 1'b1;
pika_color[9955] <= 1'b1;
pika_color[9968] <= 1'b1;
pika_color[10026] <= 1'b1;
pika_color[10030] <= 1'b1;
pika_color[10031] <= 1'b1;
pika_color[10050] <= 1'b1;
pika_color[10051] <= 1'b1;
pika_color[10054] <= 1'b1;
pika_color[10055] <= 1'b1;
pika_color[10069] <= 1'b1;
pika_color[10070] <= 1'b1;
pika_color[10083] <= 1'b1;
pika_color[10142] <= 1'b1;
pika_color[10146] <= 1'b1;
pika_color[10147] <= 1'b1;
pika_color[10167] <= 1'b1;
pika_color[10168] <= 1'b1;
pika_color[10184] <= 1'b1;
pika_color[10198] <= 1'b1;
pika_color[10257] <= 1'b1;
pika_color[10263] <= 1'b1;
pika_color[10298] <= 1'b1;
pika_color[10299] <= 1'b1;
pika_color[10313] <= 1'b1;
pika_color[10371] <= 1'b1;
pika_color[10379] <= 1'b1;
pika_color[10380] <= 1'b1;
pika_color[10381] <= 1'b1;
pika_color[10413] <= 1'b1;
pika_color[10427] <= 1'b1;
pika_color[10428] <= 1'b1;
pika_color[10485] <= 1'b1;
pika_color[10486] <= 1'b1;
pika_color[10496] <= 1'b1;
pika_color[10497] <= 1'b1;
pika_color[10526] <= 1'b1;
pika_color[10527] <= 1'b1;
pika_color[10542] <= 1'b1;
pika_color[10600] <= 1'b1;
pika_color[10641] <= 1'b1;
pika_color[10657] <= 1'b1;
pika_color[10715] <= 1'b1;
pika_color[10772] <= 1'b1;
pika_color[10830] <= 1'b1;
pika_color[10887] <= 1'b1;
pika_color[10945] <= 1'b1;
pika_color[11002] <= 1'b1;
pika_color[11060] <= 1'b1;
pika_color[11117] <= 1'b1;
pika_color[11175] <= 1'b1;
pika_color[11232] <= 1'b1;
pika_color[11290] <= 1'b1;
pika_color[11347] <= 1'b1;
pika_color[11405] <= 1'b1;
pika_color[11462] <= 1'b1;
pika_color[11520] <= 1'b1;
pika_color[11577] <= 1'b1;
pika_color[11634] <= 1'b1;
pika_color[11692] <= 1'b1;
pika_color[11748] <= 1'b1;
pika_color[11775] <= 1'b1;
pika_color[11807] <= 1'b1;
pika_color[11862] <= 1'b1;
pika_color[11863] <= 1'b1;
pika_color[11864] <= 1'b1;
pika_color[11888] <= 1'b1;
pika_color[11889] <= 1'b1;
pika_color[11890] <= 1'b1;
pika_color[11922] <= 1'b1;
pika_color[11977] <= 1'b1;
pika_color[11979] <= 1'b1;
pika_color[11980] <= 1'b1;
pika_color[12002] <= 1'b1;
pika_color[12003] <= 1'b1;
pika_color[12037] <= 1'b1;
pika_color[12092] <= 1'b1;
pika_color[12095] <= 1'b1;
pika_color[12116] <= 1'b1;
pika_color[12117] <= 1'b1;
pika_color[12152] <= 1'b1;
pika_color[12207] <= 1'b1;
pika_color[12210] <= 1'b1;
pika_color[12230] <= 1'b1;
pika_color[12231] <= 1'b1;
pika_color[12267] <= 1'b1;
pika_color[12322] <= 1'b1;
pika_color[12325] <= 1'b1;
pika_color[12344] <= 1'b1;
pika_color[12345] <= 1'b1;
pika_color[12382] <= 1'b1;
pika_color[12436] <= 1'b1;
pika_color[12437] <= 1'b1;
pika_color[12440] <= 1'b1;
pika_color[12458] <= 1'b1;
pika_color[12459] <= 1'b1;
pika_color[12497] <= 1'b1;
pika_color[12498] <= 1'b1;
pika_color[12551] <= 1'b1;
pika_color[12555] <= 1'b1;
pika_color[12556] <= 1'b1;
pika_color[12573] <= 1'b1;
pika_color[12613] <= 1'b1;
pika_color[12666] <= 1'b1;
pika_color[12671] <= 1'b1;
pika_color[12688] <= 1'b1;
pika_color[12728] <= 1'b1;
pika_color[12780] <= 1'b1;
pika_color[12781] <= 1'b1;
pika_color[12786] <= 1'b1;
pika_color[12787] <= 1'b1;
pika_color[12803] <= 1'b1;
pika_color[12843] <= 1'b1;
pika_color[12895] <= 1'b1;
pika_color[12902] <= 1'b1;
pika_color[12918] <= 1'b1;
pika_color[12958] <= 1'b1;
pika_color[13009] <= 1'b1;
pika_color[13010] <= 1'b1;
pika_color[13017] <= 1'b1;
pika_color[13033] <= 1'b1;
pika_color[13073] <= 1'b1;
pika_color[13124] <= 1'b1;
pika_color[13132] <= 1'b1;
pika_color[13148] <= 1'b1;
pika_color[13149] <= 1'b1;
pika_color[13188] <= 1'b1;
pika_color[13239] <= 1'b1;
pika_color[13247] <= 1'b1;
pika_color[13264] <= 1'b1;
pika_color[13303] <= 1'b1;
pika_color[13354] <= 1'b1;
pika_color[13362] <= 1'b1;
pika_color[13363] <= 1'b1;
pika_color[13379] <= 1'b1;
pika_color[13418] <= 1'b1;
pika_color[13469] <= 1'b1;
pika_color[13478] <= 1'b1;
pika_color[13494] <= 1'b1;
pika_color[13533] <= 1'b1;
pika_color[13583] <= 1'b1;
pika_color[13584] <= 1'b1;
pika_color[13593] <= 1'b1;
pika_color[13594] <= 1'b1;
pika_color[13609] <= 1'b1;
pika_color[13648] <= 1'b1;
pika_color[13698] <= 1'b1;
pika_color[13709] <= 1'b1;
pika_color[13724] <= 1'b1;
pika_color[13763] <= 1'b1;
pika_color[13813] <= 1'b1;
pika_color[13824] <= 1'b1;
pika_color[13839] <= 1'b1;
pika_color[13878] <= 1'b1;
pika_color[13928] <= 1'b1;
pika_color[13939] <= 1'b1;
pika_color[13940] <= 1'b1;
pika_color[13953] <= 1'b1;
pika_color[13954] <= 1'b1;
pika_color[13993] <= 1'b1;
pika_color[14043] <= 1'b1;
pika_color[14055] <= 1'b1;
pika_color[14067] <= 1'b1;
pika_color[14068] <= 1'b1;
pika_color[14108] <= 1'b1;
pika_color[14158] <= 1'b1;
pika_color[14171] <= 1'b1;
pika_color[14182] <= 1'b1;
pika_color[14223] <= 1'b1;
pika_color[14273] <= 1'b1;
pika_color[14286] <= 1'b1;
pika_color[14287] <= 1'b1;
pika_color[14295] <= 1'b1;
pika_color[14296] <= 1'b1;
pika_color[14297] <= 1'b1;
pika_color[14338] <= 1'b1;
pika_color[14388] <= 1'b1;
pika_color[14402] <= 1'b1;
pika_color[14403] <= 1'b1;
pika_color[14404] <= 1'b1;
pika_color[14405] <= 1'b1;
pika_color[14406] <= 1'b1;
pika_color[14407] <= 1'b1;
pika_color[14408] <= 1'b1;
pika_color[14409] <= 1'b1;
pika_color[14410] <= 1'b1;
pika_color[14453] <= 1'b1;
pika_color[14503] <= 1'b1;
pika_color[14522] <= 1'b1;
pika_color[14523] <= 1'b1;
pika_color[14568] <= 1'b1;
pika_color[14618] <= 1'b1;
pika_color[14619] <= 1'b1;
pika_color[14683] <= 1'b1;
pika_color[14734] <= 1'b1;
pika_color[14735] <= 1'b1;
pika_color[14798] <= 1'b1;
pika_color[14850] <= 1'b1;
pika_color[14912] <= 1'b1;
pika_color[14913] <= 1'b1;
pika_color[14965] <= 1'b1;
pika_color[14966] <= 1'b1;
pika_color[15027] <= 1'b1;
pika_color[15081] <= 1'b1;
pika_color[15082] <= 1'b1;
pika_color[15141] <= 1'b1;
pika_color[15142] <= 1'b1;
pika_color[15197] <= 1'b1;
pika_color[15198] <= 1'b1;
pika_color[15256] <= 1'b1;
pika_color[15313] <= 1'b1;
pika_color[15314] <= 1'b1;
pika_color[15370] <= 1'b1;
pika_color[15371] <= 1'b1;
pika_color[15429] <= 1'b1;
pika_color[15430] <= 1'b1;
pika_color[15431] <= 1'b1;
pika_color[15432] <= 1'b1;
pika_color[15433] <= 1'b1;
pika_color[15485] <= 1'b1;
pika_color[15548] <= 1'b1;
pika_color[15549] <= 1'b1;
pika_color[15550] <= 1'b1;
pika_color[15600] <= 1'b1;
pika_color[15665] <= 1'b1;
pika_color[15670] <= 1'b1;
pika_color[15671] <= 1'b1;
pika_color[15672] <= 1'b1;
pika_color[15673] <= 1'b1;
pika_color[15674] <= 1'b1;
pika_color[15675] <= 1'b1;
pika_color[15676] <= 1'b1;
pika_color[15677] <= 1'b1;
pika_color[15678] <= 1'b1;
pika_color[15679] <= 1'b1;
pika_color[15715] <= 1'b1;
pika_color[15780] <= 1'b1;
pika_color[15781] <= 1'b1;
pika_color[15782] <= 1'b1;
pika_color[15783] <= 1'b1;
pika_color[15784] <= 1'b1;
pika_color[15785] <= 1'b1;
pika_color[15794] <= 1'b1;
pika_color[15795] <= 1'b1;
pika_color[15796] <= 1'b1;
pika_color[15797] <= 1'b1;
pika_color[15829] <= 1'b1;
pika_color[15830] <= 1'b1;
pika_color[15912] <= 1'b1;
pika_color[15913] <= 1'b1;
pika_color[15914] <= 1'b1;
pika_color[15915] <= 1'b1;
pika_color[15916] <= 1'b1;
pika_color[15917] <= 1'b1;
pika_color[15918] <= 1'b1;
pika_color[15919] <= 1'b1;
pika_color[15943] <= 1'b1;
pika_color[16033] <= 1'b1;
pika_color[16034] <= 1'b1;
pika_color[16035] <= 1'b1;
pika_color[16036] <= 1'b1;
pika_color[16037] <= 1'b1;
pika_color[16038] <= 1'b1;
pika_color[16039] <= 1'b1;
pika_color[16057] <= 1'b1;
pika_color[16058] <= 1'b1;
pika_color[16154] <= 1'b1;
pika_color[16155] <= 1'b1;
pika_color[16156] <= 1'b1;
pika_color[16157] <= 1'b1;
pika_color[16158] <= 1'b1;
pika_color[16171] <= 1'b1;
pika_color[16172] <= 1'b1;
pika_color[16273] <= 1'b1;
pika_color[16284] <= 1'b1;
pika_color[16285] <= 1'b1;
pika_color[16286] <= 1'b1;
pika_color[16388] <= 1'b1;
pika_color[16397] <= 1'b1;
pika_color[16398] <= 1'b1;
pika_color[16399] <= 1'b1;
pika_color[16503] <= 1'b1;
pika_color[16512] <= 1'b1;
pika_color[16618] <= 1'b1;
pika_color[16627] <= 1'b1;
pika_color[16733] <= 1'b1;
pika_color[16742] <= 1'b1;
pika_color[16848] <= 1'b1;
pika_color[16849] <= 1'b1;
pika_color[16850] <= 1'b1;
pika_color[16851] <= 1'b1;
pika_color[16852] <= 1'b1;
pika_color[16853] <= 1'b1;
pika_color[16854] <= 1'b1;
pika_color[16855] <= 1'b1;
pika_color[16856] <= 1'b1;

		end
		move30, move31, move32, move33, move34, move35, move36, move37, move38, move39:
		begin
		pika_color[884] <= 1'b1;
pika_color[885] <= 1'b1;
pika_color[886] <= 1'b1;
pika_color[887] <= 1'b1;
pika_color[888] <= 1'b1;
pika_color[996] <= 1'b1;
pika_color[997] <= 1'b1;
pika_color[998] <= 1'b1;
pika_color[999] <= 1'b1;
pika_color[1000] <= 1'b1;
pika_color[1001] <= 1'b1;
pika_color[1002] <= 1'b1;
pika_color[1003] <= 1'b1;
pika_color[1004] <= 1'b1;
pika_color[1109] <= 1'b1;
pika_color[1110] <= 1'b1;
pika_color[1111] <= 1'b1;
pika_color[1112] <= 1'b1;
pika_color[1113] <= 1'b1;
pika_color[1114] <= 1'b1;
pika_color[1115] <= 1'b1;
pika_color[1116] <= 1'b1;
pika_color[1117] <= 1'b1;
pika_color[1118] <= 1'b1;
pika_color[1119] <= 1'b1;
pika_color[1120] <= 1'b1;
pika_color[1224] <= 1'b1;
pika_color[1225] <= 1'b1;
pika_color[1227] <= 1'b1;
pika_color[1228] <= 1'b1;
pika_color[1229] <= 1'b1;
pika_color[1230] <= 1'b1;
pika_color[1231] <= 1'b1;
pika_color[1232] <= 1'b1;
pika_color[1233] <= 1'b1;
pika_color[1234] <= 1'b1;
pika_color[1235] <= 1'b1;
pika_color[1338] <= 1'b1;
pika_color[1339] <= 1'b1;
pika_color[1342] <= 1'b1;
pika_color[1343] <= 1'b1;
pika_color[1344] <= 1'b1;
pika_color[1345] <= 1'b1;
pika_color[1346] <= 1'b1;
pika_color[1347] <= 1'b1;
pika_color[1348] <= 1'b1;
pika_color[1349] <= 1'b1;
pika_color[1350] <= 1'b1;
pika_color[1451] <= 1'b1;
pika_color[1452] <= 1'b1;
pika_color[1453] <= 1'b1;
pika_color[1457] <= 1'b1;
pika_color[1458] <= 1'b1;
pika_color[1459] <= 1'b1;
pika_color[1460] <= 1'b1;
pika_color[1461] <= 1'b1;
pika_color[1462] <= 1'b1;
pika_color[1463] <= 1'b1;
pika_color[1464] <= 1'b1;
pika_color[1565] <= 1'b1;
pika_color[1566] <= 1'b1;
pika_color[1572] <= 1'b1;
pika_color[1573] <= 1'b1;
pika_color[1574] <= 1'b1;
pika_color[1575] <= 1'b1;
pika_color[1576] <= 1'b1;
pika_color[1577] <= 1'b1;
pika_color[1578] <= 1'b1;
pika_color[1579] <= 1'b1;
pika_color[1679] <= 1'b1;
pika_color[1680] <= 1'b1;
pika_color[1688] <= 1'b1;
pika_color[1689] <= 1'b1;
pika_color[1690] <= 1'b1;
pika_color[1691] <= 1'b1;
pika_color[1692] <= 1'b1;
pika_color[1693] <= 1'b1;
pika_color[1694] <= 1'b1;
pika_color[1735] <= 1'b1;
pika_color[1736] <= 1'b1;
pika_color[1794] <= 1'b1;
pika_color[1803] <= 1'b1;
pika_color[1804] <= 1'b1;
pika_color[1805] <= 1'b1;
pika_color[1806] <= 1'b1;
pika_color[1807] <= 1'b1;
pika_color[1808] <= 1'b1;
pika_color[1849] <= 1'b1;
pika_color[1850] <= 1'b1;
pika_color[1851] <= 1'b1;
pika_color[1852] <= 1'b1;
pika_color[1853] <= 1'b1;
pika_color[1854] <= 1'b1;
pika_color[1908] <= 1'b1;
pika_color[1909] <= 1'b1;
pika_color[1918] <= 1'b1;
pika_color[1919] <= 1'b1;
pika_color[1920] <= 1'b1;
pika_color[1921] <= 1'b1;
pika_color[1922] <= 1'b1;
pika_color[1923] <= 1'b1;
pika_color[1964] <= 1'b1;
pika_color[1965] <= 1'b1;
pika_color[1966] <= 1'b1;
pika_color[1967] <= 1'b1;
pika_color[1968] <= 1'b1;
pika_color[1969] <= 1'b1;
pika_color[1970] <= 1'b1;
pika_color[1971] <= 1'b1;
pika_color[1972] <= 1'b1;
pika_color[2022] <= 1'b1;
pika_color[2023] <= 1'b1;
pika_color[2033] <= 1'b1;
pika_color[2034] <= 1'b1;
pika_color[2035] <= 1'b1;
pika_color[2036] <= 1'b1;
pika_color[2037] <= 1'b1;
pika_color[2079] <= 1'b1;
pika_color[2080] <= 1'b1;
pika_color[2081] <= 1'b1;
pika_color[2082] <= 1'b1;
pika_color[2083] <= 1'b1;
pika_color[2084] <= 1'b1;
pika_color[2085] <= 1'b1;
pika_color[2086] <= 1'b1;
pika_color[2087] <= 1'b1;
pika_color[2088] <= 1'b1;
pika_color[2136] <= 1'b1;
pika_color[2137] <= 1'b1;
pika_color[2148] <= 1'b1;
pika_color[2149] <= 1'b1;
pika_color[2150] <= 1'b1;
pika_color[2151] <= 1'b1;
pika_color[2152] <= 1'b1;
pika_color[2194] <= 1'b1;
pika_color[2195] <= 1'b1;
pika_color[2196] <= 1'b1;
pika_color[2197] <= 1'b1;
pika_color[2198] <= 1'b1;
pika_color[2199] <= 1'b1;
pika_color[2200] <= 1'b1;
pika_color[2203] <= 1'b1;
pika_color[2204] <= 1'b1;
pika_color[2205] <= 1'b1;
pika_color[2251] <= 1'b1;
pika_color[2263] <= 1'b1;
pika_color[2264] <= 1'b1;
pika_color[2265] <= 1'b1;
pika_color[2266] <= 1'b1;
pika_color[2267] <= 1'b1;
pika_color[2309] <= 1'b1;
pika_color[2310] <= 1'b1;
pika_color[2311] <= 1'b1;
pika_color[2312] <= 1'b1;
pika_color[2313] <= 1'b1;
pika_color[2314] <= 1'b1;
pika_color[2315] <= 1'b1;
pika_color[2319] <= 1'b1;
pika_color[2320] <= 1'b1;
pika_color[2321] <= 1'b1;
pika_color[2365] <= 1'b1;
pika_color[2379] <= 1'b1;
pika_color[2380] <= 1'b1;
pika_color[2381] <= 1'b1;
pika_color[2424] <= 1'b1;
pika_color[2425] <= 1'b1;
pika_color[2426] <= 1'b1;
pika_color[2427] <= 1'b1;
pika_color[2428] <= 1'b1;
pika_color[2429] <= 1'b1;
pika_color[2436] <= 1'b1;
pika_color[2437] <= 1'b1;
pika_color[2480] <= 1'b1;
pika_color[2494] <= 1'b1;
pika_color[2495] <= 1'b1;
pika_color[2496] <= 1'b1;
pika_color[2539] <= 1'b1;
pika_color[2540] <= 1'b1;
pika_color[2541] <= 1'b1;
pika_color[2542] <= 1'b1;
pika_color[2543] <= 1'b1;
pika_color[2544] <= 1'b1;
pika_color[2552] <= 1'b1;
pika_color[2553] <= 1'b1;
pika_color[2594] <= 1'b1;
pika_color[2595] <= 1'b1;
pika_color[2610] <= 1'b1;
pika_color[2611] <= 1'b1;
pika_color[2655] <= 1'b1;
pika_color[2656] <= 1'b1;
pika_color[2657] <= 1'b1;
pika_color[2658] <= 1'b1;
pika_color[2668] <= 1'b1;
pika_color[2709] <= 1'b1;
pika_color[2724] <= 1'b1;
pika_color[2725] <= 1'b1;
pika_color[2770] <= 1'b1;
pika_color[2771] <= 1'b1;
pika_color[2772] <= 1'b1;
pika_color[2773] <= 1'b1;
pika_color[2783] <= 1'b1;
pika_color[2784] <= 1'b1;
pika_color[2823] <= 1'b1;
pika_color[2824] <= 1'b1;
pika_color[2839] <= 1'b1;
pika_color[2840] <= 1'b1;
pika_color[2885] <= 1'b1;
pika_color[2886] <= 1'b1;
pika_color[2887] <= 1'b1;
pika_color[2888] <= 1'b1;
pika_color[2899] <= 1'b1;
pika_color[2938] <= 1'b1;
pika_color[2954] <= 1'b1;
pika_color[3000] <= 1'b1;
pika_color[3001] <= 1'b1;
pika_color[3002] <= 1'b1;
pika_color[3003] <= 1'b1;
pika_color[3014] <= 1'b1;
pika_color[3015] <= 1'b1;
pika_color[3052] <= 1'b1;
pika_color[3053] <= 1'b1;
pika_color[3068] <= 1'b1;
pika_color[3069] <= 1'b1;
pika_color[3116] <= 1'b1;
pika_color[3117] <= 1'b1;
pika_color[3118] <= 1'b1;
pika_color[3130] <= 1'b1;
pika_color[3167] <= 1'b1;
pika_color[3183] <= 1'b1;
pika_color[3231] <= 1'b1;
pika_color[3232] <= 1'b1;
pika_color[3245] <= 1'b1;
pika_color[3246] <= 1'b1;
pika_color[3281] <= 1'b1;
pika_color[3297] <= 1'b1;
pika_color[3346] <= 1'b1;
pika_color[3347] <= 1'b1;
pika_color[3361] <= 1'b1;
pika_color[3362] <= 1'b1;
pika_color[3396] <= 1'b1;
pika_color[3411] <= 1'b1;
pika_color[3412] <= 1'b1;
pika_color[3462] <= 1'b1;
pika_color[3477] <= 1'b1;
pika_color[3478] <= 1'b1;
pika_color[3510] <= 1'b1;
pika_color[3511] <= 1'b1;
pika_color[3525] <= 1'b1;
pika_color[3526] <= 1'b1;
pika_color[3577] <= 1'b1;
pika_color[3578] <= 1'b1;
pika_color[3593] <= 1'b1;
pika_color[3608] <= 1'b1;
pika_color[3609] <= 1'b1;
pika_color[3610] <= 1'b1;
pika_color[3611] <= 1'b1;
pika_color[3612] <= 1'b1;
pika_color[3613] <= 1'b1;
pika_color[3614] <= 1'b1;
pika_color[3615] <= 1'b1;
pika_color[3616] <= 1'b1;
pika_color[3617] <= 1'b1;
pika_color[3625] <= 1'b1;
pika_color[3640] <= 1'b1;
pika_color[3693] <= 1'b1;
pika_color[3694] <= 1'b1;
pika_color[3708] <= 1'b1;
pika_color[3709] <= 1'b1;
pika_color[3721] <= 1'b1;
pika_color[3722] <= 1'b1;
pika_color[3723] <= 1'b1;
pika_color[3732] <= 1'b1;
pika_color[3733] <= 1'b1;
pika_color[3734] <= 1'b1;
pika_color[3735] <= 1'b1;
pika_color[3740] <= 1'b1;
pika_color[3754] <= 1'b1;
pika_color[3809] <= 1'b1;
pika_color[3824] <= 1'b1;
pika_color[3833] <= 1'b1;
pika_color[3834] <= 1'b1;
pika_color[3835] <= 1'b1;
pika_color[3836] <= 1'b1;
pika_color[3850] <= 1'b1;
pika_color[3851] <= 1'b1;
pika_color[3852] <= 1'b1;
pika_color[3855] <= 1'b1;
pika_color[3868] <= 1'b1;
pika_color[3869] <= 1'b1;
pika_color[3924] <= 1'b1;
pika_color[3925] <= 1'b1;
pika_color[3939] <= 1'b1;
pika_color[3940] <= 1'b1;
pika_color[3945] <= 1'b1;
pika_color[3946] <= 1'b1;
pika_color[3947] <= 1'b1;
pika_color[3948] <= 1'b1;
pika_color[3967] <= 1'b1;
pika_color[3968] <= 1'b1;
pika_color[3969] <= 1'b1;
pika_color[3970] <= 1'b1;
pika_color[3983] <= 1'b1;
pika_color[4040] <= 1'b1;
pika_color[4055] <= 1'b1;
pika_color[4056] <= 1'b1;
pika_color[4058] <= 1'b1;
pika_color[4059] <= 1'b1;
pika_color[4060] <= 1'b1;
pika_color[4085] <= 1'b1;
pika_color[4097] <= 1'b1;
pika_color[4098] <= 1'b1;
pika_color[4155] <= 1'b1;
pika_color[4156] <= 1'b1;
pika_color[4171] <= 1'b1;
pika_color[4172] <= 1'b1;
pika_color[4173] <= 1'b1;
pika_color[4212] <= 1'b1;
pika_color[4271] <= 1'b1;
pika_color[4286] <= 1'b1;
pika_color[4287] <= 1'b1;
pika_color[4326] <= 1'b1;
pika_color[4327] <= 1'b1;
pika_color[4386] <= 1'b1;
pika_color[4387] <= 1'b1;
pika_color[4402] <= 1'b1;
pika_color[4403] <= 1'b1;
pika_color[4440] <= 1'b1;
pika_color[4502] <= 1'b1;
pika_color[4503] <= 1'b1;
pika_color[4518] <= 1'b1;
pika_color[4554] <= 1'b1;
pika_color[4555] <= 1'b1;
pika_color[4617] <= 1'b1;
pika_color[4618] <= 1'b1;
pika_color[4619] <= 1'b1;
pika_color[4633] <= 1'b1;
pika_color[4668] <= 1'b1;
pika_color[4669] <= 1'b1;
pika_color[4732] <= 1'b1;
pika_color[4734] <= 1'b1;
pika_color[4783] <= 1'b1;
pika_color[4784] <= 1'b1;
pika_color[4847] <= 1'b1;
pika_color[4849] <= 1'b1;
pika_color[4850] <= 1'b1;
pika_color[4899] <= 1'b1;
pika_color[4900] <= 1'b1;
pika_color[4962] <= 1'b1;
pika_color[4965] <= 1'b1;
pika_color[4966] <= 1'b1;
pika_color[5015] <= 1'b1;
pika_color[5016] <= 1'b1;
pika_color[5077] <= 1'b1;
pika_color[5078] <= 1'b1;
pika_color[5081] <= 1'b1;
pika_color[5082] <= 1'b1;
pika_color[5083] <= 1'b1;
pika_color[5131] <= 1'b1;
pika_color[5193] <= 1'b1;
pika_color[5198] <= 1'b1;
pika_color[5199] <= 1'b1;
pika_color[5246] <= 1'b1;
pika_color[5247] <= 1'b1;
pika_color[5308] <= 1'b1;
pika_color[5314] <= 1'b1;
pika_color[5362] <= 1'b1;
pika_color[5423] <= 1'b1;
pika_color[5424] <= 1'b1;
pika_color[5430] <= 1'b1;
pika_color[5477] <= 1'b1;
pika_color[5539] <= 1'b1;
pika_color[5545] <= 1'b1;
pika_color[5592] <= 1'b1;
pika_color[5593] <= 1'b1;
pika_color[5654] <= 1'b1;
pika_color[5659] <= 1'b1;
pika_color[5708] <= 1'b1;
pika_color[5769] <= 1'b1;
pika_color[5770] <= 1'b1;
pika_color[5774] <= 1'b1;
pika_color[5823] <= 1'b1;
pika_color[5824] <= 1'b1;
pika_color[5885] <= 1'b1;
pika_color[5889] <= 1'b1;
pika_color[5939] <= 1'b1;
pika_color[6000] <= 1'b1;
pika_color[6004] <= 1'b1;
pika_color[6054] <= 1'b1;
pika_color[6115] <= 1'b1;
pika_color[6119] <= 1'b1;
pika_color[6169] <= 1'b1;
pika_color[6170] <= 1'b1;
pika_color[6230] <= 1'b1;
pika_color[6234] <= 1'b1;
pika_color[6285] <= 1'b1;
pika_color[6345] <= 1'b1;
pika_color[6349] <= 1'b1;
pika_color[6386] <= 1'b1;
pika_color[6387] <= 1'b1;
pika_color[6388] <= 1'b1;
pika_color[6399] <= 1'b1;
pika_color[6400] <= 1'b1;
pika_color[6460] <= 1'b1;
pika_color[6461] <= 1'b1;
pika_color[6464] <= 1'b1;
pika_color[6499] <= 1'b1;
pika_color[6500] <= 1'b1;
pika_color[6501] <= 1'b1;
pika_color[6502] <= 1'b1;
pika_color[6503] <= 1'b1;
pika_color[6510] <= 1'b1;
pika_color[6511] <= 1'b1;
pika_color[6512] <= 1'b1;
pika_color[6513] <= 1'b1;
pika_color[6514] <= 1'b1;
pika_color[6515] <= 1'b1;
pika_color[6516] <= 1'b1;
pika_color[6517] <= 1'b1;
pika_color[6518] <= 1'b1;
pika_color[6576] <= 1'b1;
pika_color[6579] <= 1'b1;
pika_color[6613] <= 1'b1;
pika_color[6614] <= 1'b1;
pika_color[6615] <= 1'b1;
pika_color[6624] <= 1'b1;
pika_color[6625] <= 1'b1;
pika_color[6633] <= 1'b1;
pika_color[6634] <= 1'b1;
pika_color[6691] <= 1'b1;
pika_color[6694] <= 1'b1;
pika_color[6738] <= 1'b1;
pika_color[6739] <= 1'b1;
pika_color[6749] <= 1'b1;
pika_color[6750] <= 1'b1;
pika_color[6806] <= 1'b1;
pika_color[6807] <= 1'b1;
pika_color[6809] <= 1'b1;
pika_color[6810] <= 1'b1;
pika_color[6852] <= 1'b1;
pika_color[6853] <= 1'b1;
pika_color[6865] <= 1'b1;
pika_color[6922] <= 1'b1;
pika_color[6925] <= 1'b1;
pika_color[6967] <= 1'b1;
pika_color[6980] <= 1'b1;
pika_color[6981] <= 1'b1;
pika_color[7037] <= 1'b1;
pika_color[7040] <= 1'b1;
pika_color[7052] <= 1'b1;
pika_color[7053] <= 1'b1;
pika_color[7054] <= 1'b1;
pika_color[7055] <= 1'b1;
pika_color[7056] <= 1'b1;
pika_color[7082] <= 1'b1;
pika_color[7096] <= 1'b1;
pika_color[7097] <= 1'b1;
pika_color[7152] <= 1'b1;
pika_color[7153] <= 1'b1;
pika_color[7155] <= 1'b1;
pika_color[7164] <= 1'b1;
pika_color[7165] <= 1'b1;
pika_color[7166] <= 1'b1;
pika_color[7167] <= 1'b1;
pika_color[7168] <= 1'b1;
pika_color[7169] <= 1'b1;
pika_color[7170] <= 1'b1;
pika_color[7171] <= 1'b1;
pika_color[7197] <= 1'b1;
pika_color[7198] <= 1'b1;
pika_color[7212] <= 1'b1;
pika_color[7268] <= 1'b1;
pika_color[7270] <= 1'b1;
pika_color[7293] <= 1'b1;
pika_color[7294] <= 1'b1;
pika_color[7295] <= 1'b1;
pika_color[7296] <= 1'b1;
pika_color[7313] <= 1'b1;
pika_color[7327] <= 1'b1;
pika_color[7383] <= 1'b1;
pika_color[7385] <= 1'b1;
pika_color[7407] <= 1'b1;
pika_color[7408] <= 1'b1;
pika_color[7409] <= 1'b1;
pika_color[7410] <= 1'b1;
pika_color[7411] <= 1'b1;
pika_color[7428] <= 1'b1;
pika_color[7442] <= 1'b1;
pika_color[7443] <= 1'b1;
pika_color[7498] <= 1'b1;
pika_color[7500] <= 1'b1;
pika_color[7524] <= 1'b1;
pika_color[7525] <= 1'b1;
pika_color[7543] <= 1'b1;
pika_color[7544] <= 1'b1;
pika_color[7558] <= 1'b1;
pika_color[7613] <= 1'b1;
pika_color[7614] <= 1'b1;
pika_color[7615] <= 1'b1;
pika_color[7659] <= 1'b1;
pika_color[7673] <= 1'b1;
pika_color[7729] <= 1'b1;
pika_color[7730] <= 1'b1;
pika_color[7731] <= 1'b1;
pika_color[7774] <= 1'b1;
pika_color[7788] <= 1'b1;
pika_color[7845] <= 1'b1;
pika_color[7846] <= 1'b1;
pika_color[7872] <= 1'b1;
pika_color[7873] <= 1'b1;
pika_color[7874] <= 1'b1;
pika_color[7875] <= 1'b1;
pika_color[7889] <= 1'b1;
pika_color[7890] <= 1'b1;
pika_color[7903] <= 1'b1;
pika_color[7961] <= 1'b1;
pika_color[7984] <= 1'b1;
pika_color[7985] <= 1'b1;
pika_color[7986] <= 1'b1;
pika_color[7990] <= 1'b1;
pika_color[7991] <= 1'b1;
pika_color[7992] <= 1'b1;
pika_color[8005] <= 1'b1;
pika_color[8018] <= 1'b1;
pika_color[8076] <= 1'b1;
pika_color[8098] <= 1'b1;
pika_color[8099] <= 1'b1;
pika_color[8107] <= 1'b1;
pika_color[8120] <= 1'b1;
pika_color[8133] <= 1'b1;
pika_color[8191] <= 1'b1;
pika_color[8210] <= 1'b1;
pika_color[8211] <= 1'b1;
pika_color[8212] <= 1'b1;
pika_color[8216] <= 1'b1;
pika_color[8217] <= 1'b1;
pika_color[8218] <= 1'b1;
pika_color[8219] <= 1'b1;
pika_color[8222] <= 1'b1;
pika_color[8235] <= 1'b1;
pika_color[8248] <= 1'b1;
pika_color[8306] <= 1'b1;
pika_color[8307] <= 1'b1;
pika_color[8325] <= 1'b1;
pika_color[8329] <= 1'b1;
pika_color[8330] <= 1'b1;
pika_color[8335] <= 1'b1;
pika_color[8336] <= 1'b1;
pika_color[8349] <= 1'b1;
pika_color[8350] <= 1'b1;
pika_color[8363] <= 1'b1;
pika_color[8422] <= 1'b1;
pika_color[8441] <= 1'b1;
pika_color[8442] <= 1'b1;
pika_color[8443] <= 1'b1;
pika_color[8444] <= 1'b1;
pika_color[8450] <= 1'b1;
pika_color[8464] <= 1'b1;
pika_color[8478] <= 1'b1;
pika_color[8537] <= 1'b1;
pika_color[8558] <= 1'b1;
pika_color[8559] <= 1'b1;
pika_color[8564] <= 1'b1;
pika_color[8579] <= 1'b1;
pika_color[8593] <= 1'b1;
pika_color[8652] <= 1'b1;
pika_color[8653] <= 1'b1;
pika_color[8675] <= 1'b1;
pika_color[8676] <= 1'b1;
pika_color[8677] <= 1'b1;
pika_color[8678] <= 1'b1;
pika_color[8693] <= 1'b1;
pika_color[8694] <= 1'b1;
pika_color[8708] <= 1'b1;
pika_color[8709] <= 1'b1;
pika_color[8768] <= 1'b1;
pika_color[8808] <= 1'b1;
pika_color[8824] <= 1'b1;
pika_color[8883] <= 1'b1;
pika_color[8884] <= 1'b1;
pika_color[8922] <= 1'b1;
pika_color[8923] <= 1'b1;
pika_color[8939] <= 1'b1;
pika_color[8999] <= 1'b1;
pika_color[9000] <= 1'b1;
pika_color[9001] <= 1'b1;
pika_color[9037] <= 1'b1;
pika_color[9054] <= 1'b1;
pika_color[9115] <= 1'b1;
pika_color[9116] <= 1'b1;
pika_color[9117] <= 1'b1;
pika_color[9151] <= 1'b1;
pika_color[9152] <= 1'b1;
pika_color[9169] <= 1'b1;
pika_color[9230] <= 1'b1;
pika_color[9232] <= 1'b1;
pika_color[9233] <= 1'b1;
pika_color[9265] <= 1'b1;
pika_color[9266] <= 1'b1;
pika_color[9284] <= 1'b1;
pika_color[9344] <= 1'b1;
pika_color[9348] <= 1'b1;
pika_color[9349] <= 1'b1;
pika_color[9350] <= 1'b1;
pika_color[9351] <= 1'b1;
pika_color[9380] <= 1'b1;
pika_color[9399] <= 1'b1;
pika_color[9459] <= 1'b1;
pika_color[9466] <= 1'b1;
pika_color[9467] <= 1'b1;
pika_color[9514] <= 1'b1;
pika_color[9574] <= 1'b1;
pika_color[9629] <= 1'b1;
pika_color[9688] <= 1'b1;
pika_color[9689] <= 1'b1;
pika_color[9744] <= 1'b1;
pika_color[9745] <= 1'b1;
pika_color[9803] <= 1'b1;
pika_color[9860] <= 1'b1;
pika_color[9918] <= 1'b1;
pika_color[9975] <= 1'b1;
pika_color[10032] <= 1'b1;
pika_color[10033] <= 1'b1;
pika_color[10090] <= 1'b1;
pika_color[10147] <= 1'b1;
pika_color[10205] <= 1'b1;
pika_color[10206] <= 1'b1;
pika_color[10262] <= 1'b1;
pika_color[10321] <= 1'b1;
pika_color[10377] <= 1'b1;
pika_color[10436] <= 1'b1;
pika_color[10492] <= 1'b1;
pika_color[10512] <= 1'b1;
pika_color[10551] <= 1'b1;
pika_color[10607] <= 1'b1;
pika_color[10626] <= 1'b1;
pika_color[10627] <= 1'b1;
pika_color[10666] <= 1'b1;
pika_color[10667] <= 1'b1;
pika_color[10722] <= 1'b1;
pika_color[10741] <= 1'b1;
pika_color[10782] <= 1'b1;
pika_color[10837] <= 1'b1;
pika_color[10838] <= 1'b1;
pika_color[10855] <= 1'b1;
pika_color[10897] <= 1'b1;
pika_color[10953] <= 1'b1;
pika_color[10970] <= 1'b1;
pika_color[11012] <= 1'b1;
pika_color[11068] <= 1'b1;
pika_color[11085] <= 1'b1;
pika_color[11127] <= 1'b1;
pika_color[11183] <= 1'b1;
pika_color[11200] <= 1'b1;
pika_color[11242] <= 1'b1;
pika_color[11298] <= 1'b1;
pika_color[11315] <= 1'b1;
pika_color[11357] <= 1'b1;
pika_color[11413] <= 1'b1;
pika_color[11430] <= 1'b1;
pika_color[11472] <= 1'b1;
pika_color[11528] <= 1'b1;
pika_color[11545] <= 1'b1;
pika_color[11587] <= 1'b1;
pika_color[11588] <= 1'b1;
pika_color[11643] <= 1'b1;
pika_color[11644] <= 1'b1;
pika_color[11660] <= 1'b1;
pika_color[11703] <= 1'b1;
pika_color[11757] <= 1'b1;
pika_color[11758] <= 1'b1;
pika_color[11759] <= 1'b1;
pika_color[11775] <= 1'b1;
pika_color[11818] <= 1'b1;
pika_color[11872] <= 1'b1;
pika_color[11874] <= 1'b1;
pika_color[11890] <= 1'b1;
pika_color[11933] <= 1'b1;
pika_color[11987] <= 1'b1;
pika_color[11989] <= 1'b1;
pika_color[12005] <= 1'b1;
pika_color[12048] <= 1'b1;
pika_color[12102] <= 1'b1;
pika_color[12104] <= 1'b1;
pika_color[12105] <= 1'b1;
pika_color[12120] <= 1'b1;
pika_color[12163] <= 1'b1;
pika_color[12217] <= 1'b1;
pika_color[12220] <= 1'b1;
pika_color[12235] <= 1'b1;
pika_color[12278] <= 1'b1;
pika_color[12332] <= 1'b1;
pika_color[12335] <= 1'b1;
pika_color[12336] <= 1'b1;
pika_color[12350] <= 1'b1;
pika_color[12394] <= 1'b1;
pika_color[12447] <= 1'b1;
pika_color[12448] <= 1'b1;
pika_color[12451] <= 1'b1;
pika_color[12465] <= 1'b1;
pika_color[12509] <= 1'b1;
pika_color[12563] <= 1'b1;
pika_color[12566] <= 1'b1;
pika_color[12580] <= 1'b1;
pika_color[12624] <= 1'b1;
pika_color[12678] <= 1'b1;
pika_color[12681] <= 1'b1;
pika_color[12682] <= 1'b1;
pika_color[12694] <= 1'b1;
pika_color[12695] <= 1'b1;
pika_color[12739] <= 1'b1;
pika_color[12793] <= 1'b1;
pika_color[12797] <= 1'b1;
pika_color[12809] <= 1'b1;
pika_color[12854] <= 1'b1;
pika_color[12908] <= 1'b1;
pika_color[12912] <= 1'b1;
pika_color[12913] <= 1'b1;
pika_color[12924] <= 1'b1;
pika_color[12969] <= 1'b1;
pika_color[13023] <= 1'b1;
pika_color[13028] <= 1'b1;
pika_color[13038] <= 1'b1;
pika_color[13039] <= 1'b1;
pika_color[13084] <= 1'b1;
pika_color[13138] <= 1'b1;
pika_color[13143] <= 1'b1;
pika_color[13144] <= 1'b1;
pika_color[13152] <= 1'b1;
pika_color[13153] <= 1'b1;
pika_color[13199] <= 1'b1;
pika_color[13253] <= 1'b1;
pika_color[13254] <= 1'b1;
pika_color[13259] <= 1'b1;
pika_color[13260] <= 1'b1;
pika_color[13266] <= 1'b1;
pika_color[13267] <= 1'b1;
pika_color[13314] <= 1'b1;
pika_color[13369] <= 1'b1;
pika_color[13375] <= 1'b1;
pika_color[13376] <= 1'b1;
pika_color[13377] <= 1'b1;
pika_color[13380] <= 1'b1;
pika_color[13381] <= 1'b1;
pika_color[13429] <= 1'b1;
pika_color[13484] <= 1'b1;
pika_color[13492] <= 1'b1;
pika_color[13493] <= 1'b1;
pika_color[13494] <= 1'b1;
pika_color[13495] <= 1'b1;
pika_color[13544] <= 1'b1;
pika_color[13599] <= 1'b1;
pika_color[13659] <= 1'b1;
pika_color[13714] <= 1'b1;
pika_color[13773] <= 1'b1;
pika_color[13774] <= 1'b1;
pika_color[13829] <= 1'b1;
pika_color[13888] <= 1'b1;
pika_color[13889] <= 1'b1;
pika_color[13945] <= 1'b1;
pika_color[14003] <= 1'b1;
pika_color[14060] <= 1'b1;
pika_color[14118] <= 1'b1;
pika_color[14175] <= 1'b1;
pika_color[14232] <= 1'b1;
pika_color[14290] <= 1'b1;
pika_color[14291] <= 1'b1;
pika_color[14347] <= 1'b1;
pika_color[14406] <= 1'b1;
pika_color[14462] <= 1'b1;
pika_color[14521] <= 1'b1;
pika_color[14522] <= 1'b1;
pika_color[14577] <= 1'b1;
pika_color[14637] <= 1'b1;
pika_color[14638] <= 1'b1;
pika_color[14692] <= 1'b1;
pika_color[14753] <= 1'b1;
pika_color[14806] <= 1'b1;
pika_color[14869] <= 1'b1;
pika_color[14920] <= 1'b1;
pika_color[14921] <= 1'b1;
pika_color[14984] <= 1'b1;
pika_color[14985] <= 1'b1;
pika_color[15035] <= 1'b1;
pika_color[15100] <= 1'b1;
pika_color[15149] <= 1'b1;
pika_color[15150] <= 1'b1;
pika_color[15215] <= 1'b1;
pika_color[15216] <= 1'b1;
pika_color[15264] <= 1'b1;
pika_color[15331] <= 1'b1;
pika_color[15332] <= 1'b1;
pika_color[15333] <= 1'b1;
pika_color[15334] <= 1'b1;
pika_color[15335] <= 1'b1;
pika_color[15336] <= 1'b1;
pika_color[15345] <= 1'b1;
pika_color[15346] <= 1'b1;
pika_color[15347] <= 1'b1;
pika_color[15348] <= 1'b1;
pika_color[15349] <= 1'b1;
pika_color[15350] <= 1'b1;
pika_color[15351] <= 1'b1;
pika_color[15352] <= 1'b1;
pika_color[15353] <= 1'b1;
pika_color[15354] <= 1'b1;
pika_color[15355] <= 1'b1;
pika_color[15356] <= 1'b1;
pika_color[15357] <= 1'b1;
pika_color[15358] <= 1'b1;
pika_color[15359] <= 1'b1;
pika_color[15360] <= 1'b1;
pika_color[15361] <= 1'b1;
pika_color[15378] <= 1'b1;
pika_color[15379] <= 1'b1;
pika_color[15451] <= 1'b1;
pika_color[15459] <= 1'b1;
pika_color[15460] <= 1'b1;
pika_color[15476] <= 1'b1;
pika_color[15477] <= 1'b1;
pika_color[15478] <= 1'b1;
pika_color[15492] <= 1'b1;
pika_color[15493] <= 1'b1;
pika_color[15566] <= 1'b1;
pika_color[15575] <= 1'b1;
pika_color[15576] <= 1'b1;
pika_color[15594] <= 1'b1;
pika_color[15595] <= 1'b1;
pika_color[15596] <= 1'b1;
pika_color[15597] <= 1'b1;
pika_color[15605] <= 1'b1;
pika_color[15606] <= 1'b1;
pika_color[15607] <= 1'b1;
pika_color[15681] <= 1'b1;
pika_color[15691] <= 1'b1;
pika_color[15711] <= 1'b1;
pika_color[15712] <= 1'b1;
pika_color[15713] <= 1'b1;
pika_color[15714] <= 1'b1;
pika_color[15715] <= 1'b1;
pika_color[15716] <= 1'b1;
pika_color[15717] <= 1'b1;
pika_color[15718] <= 1'b1;
pika_color[15719] <= 1'b1;
pika_color[15720] <= 1'b1;
pika_color[15796] <= 1'b1;
pika_color[15797] <= 1'b1;
pika_color[15798] <= 1'b1;
pika_color[15799] <= 1'b1;
pika_color[15800] <= 1'b1;
pika_color[15801] <= 1'b1;
pika_color[15802] <= 1'b1;
pika_color[15805] <= 1'b1;
pika_color[15806] <= 1'b1;
pika_color[15917] <= 1'b1;
pika_color[15918] <= 1'b1;
pika_color[15919] <= 1'b1;
pika_color[15920] <= 1'b1;

		end
		move40, move41, move42, move43, move44, move45, move46, move47, move48, move49:
		begin
		pika_color[1589] <= 1'b1;
pika_color[1590] <= 1'b1;
pika_color[1591] <= 1'b1;
pika_color[1701] <= 1'b1;
pika_color[1702] <= 1'b1;
pika_color[1703] <= 1'b1;
pika_color[1704] <= 1'b1;
pika_color[1705] <= 1'b1;
pika_color[1706] <= 1'b1;
pika_color[1707] <= 1'b1;
pika_color[1708] <= 1'b1;
pika_color[1814] <= 1'b1;
pika_color[1815] <= 1'b1;
pika_color[1816] <= 1'b1;
pika_color[1817] <= 1'b1;
pika_color[1818] <= 1'b1;
pika_color[1819] <= 1'b1;
pika_color[1820] <= 1'b1;
pika_color[1821] <= 1'b1;
pika_color[1822] <= 1'b1;
pika_color[1823] <= 1'b1;
pika_color[1927] <= 1'b1;
pika_color[1928] <= 1'b1;
pika_color[1929] <= 1'b1;
pika_color[1931] <= 1'b1;
pika_color[1932] <= 1'b1;
pika_color[1933] <= 1'b1;
pika_color[1934] <= 1'b1;
pika_color[1935] <= 1'b1;
pika_color[1936] <= 1'b1;
pika_color[1937] <= 1'b1;
pika_color[1938] <= 1'b1;
pika_color[2041] <= 1'b1;
pika_color[2042] <= 1'b1;
pika_color[2046] <= 1'b1;
pika_color[2047] <= 1'b1;
pika_color[2048] <= 1'b1;
pika_color[2049] <= 1'b1;
pika_color[2050] <= 1'b1;
pika_color[2051] <= 1'b1;
pika_color[2052] <= 1'b1;
pika_color[2053] <= 1'b1;
pika_color[2154] <= 1'b1;
pika_color[2155] <= 1'b1;
pika_color[2156] <= 1'b1;
pika_color[2161] <= 1'b1;
pika_color[2162] <= 1'b1;
pika_color[2163] <= 1'b1;
pika_color[2164] <= 1'b1;
pika_color[2165] <= 1'b1;
pika_color[2166] <= 1'b1;
pika_color[2167] <= 1'b1;
pika_color[2168] <= 1'b1;
pika_color[2209] <= 1'b1;
pika_color[2210] <= 1'b1;
pika_color[2211] <= 1'b1;
pika_color[2212] <= 1'b1;
pika_color[2213] <= 1'b1;
pika_color[2214] <= 1'b1;
pika_color[2268] <= 1'b1;
pika_color[2269] <= 1'b1;
pika_color[2276] <= 1'b1;
pika_color[2277] <= 1'b1;
pika_color[2278] <= 1'b1;
pika_color[2279] <= 1'b1;
pika_color[2280] <= 1'b1;
pika_color[2281] <= 1'b1;
pika_color[2282] <= 1'b1;
pika_color[2323] <= 1'b1;
pika_color[2324] <= 1'b1;
pika_color[2329] <= 1'b1;
pika_color[2330] <= 1'b1;
pika_color[2381] <= 1'b1;
pika_color[2382] <= 1'b1;
pika_color[2383] <= 1'b1;
pika_color[2391] <= 1'b1;
pika_color[2392] <= 1'b1;
pika_color[2393] <= 1'b1;
pika_color[2394] <= 1'b1;
pika_color[2395] <= 1'b1;
pika_color[2396] <= 1'b1;
pika_color[2397] <= 1'b1;
pika_color[2438] <= 1'b1;
pika_color[2446] <= 1'b1;
pika_color[2495] <= 1'b1;
pika_color[2496] <= 1'b1;
pika_color[2506] <= 1'b1;
pika_color[2507] <= 1'b1;
pika_color[2508] <= 1'b1;
pika_color[2509] <= 1'b1;
pika_color[2510] <= 1'b1;
pika_color[2511] <= 1'b1;
pika_color[2553] <= 1'b1;
pika_color[2561] <= 1'b1;
pika_color[2562] <= 1'b1;
pika_color[2609] <= 1'b1;
pika_color[2610] <= 1'b1;
pika_color[2620] <= 1'b1;
pika_color[2621] <= 1'b1;
pika_color[2622] <= 1'b1;
pika_color[2623] <= 1'b1;
pika_color[2624] <= 1'b1;
pika_color[2625] <= 1'b1;
pika_color[2626] <= 1'b1;
pika_color[2668] <= 1'b1;
pika_color[2677] <= 1'b1;
pika_color[2678] <= 1'b1;
pika_color[2679] <= 1'b1;
pika_color[2723] <= 1'b1;
pika_color[2724] <= 1'b1;
pika_color[2735] <= 1'b1;
pika_color[2736] <= 1'b1;
pika_color[2737] <= 1'b1;
pika_color[2738] <= 1'b1;
pika_color[2739] <= 1'b1;
pika_color[2740] <= 1'b1;
pika_color[2741] <= 1'b1;
pika_color[2783] <= 1'b1;
pika_color[2794] <= 1'b1;
pika_color[2837] <= 1'b1;
pika_color[2838] <= 1'b1;
pika_color[2850] <= 1'b1;
pika_color[2851] <= 1'b1;
pika_color[2852] <= 1'b1;
pika_color[2853] <= 1'b1;
pika_color[2854] <= 1'b1;
pika_color[2855] <= 1'b1;
pika_color[2884] <= 1'b1;
pika_color[2885] <= 1'b1;
pika_color[2886] <= 1'b1;
pika_color[2887] <= 1'b1;
pika_color[2888] <= 1'b1;
pika_color[2889] <= 1'b1;
pika_color[2890] <= 1'b1;
pika_color[2891] <= 1'b1;
pika_color[2898] <= 1'b1;
pika_color[2909] <= 1'b1;
pika_color[2910] <= 1'b1;
pika_color[2951] <= 1'b1;
pika_color[2952] <= 1'b1;
pika_color[2965] <= 1'b1;
pika_color[2966] <= 1'b1;
pika_color[2967] <= 1'b1;
pika_color[2968] <= 1'b1;
pika_color[2969] <= 1'b1;
pika_color[2999] <= 1'b1;
pika_color[3000] <= 1'b1;
pika_color[3001] <= 1'b1;
pika_color[3002] <= 1'b1;
pika_color[3003] <= 1'b1;
pika_color[3004] <= 1'b1;
pika_color[3005] <= 1'b1;
pika_color[3006] <= 1'b1;
pika_color[3007] <= 1'b1;
pika_color[3008] <= 1'b1;
pika_color[3013] <= 1'b1;
pika_color[3025] <= 1'b1;
pika_color[3026] <= 1'b1;
pika_color[3027] <= 1'b1;
pika_color[3065] <= 1'b1;
pika_color[3066] <= 1'b1;
pika_color[3080] <= 1'b1;
pika_color[3081] <= 1'b1;
pika_color[3082] <= 1'b1;
pika_color[3083] <= 1'b1;
pika_color[3084] <= 1'b1;
pika_color[3114] <= 1'b1;
pika_color[3115] <= 1'b1;
pika_color[3116] <= 1'b1;
pika_color[3117] <= 1'b1;
pika_color[3118] <= 1'b1;
pika_color[3119] <= 1'b1;
pika_color[3120] <= 1'b1;
pika_color[3123] <= 1'b1;
pika_color[3124] <= 1'b1;
pika_color[3125] <= 1'b1;
pika_color[3128] <= 1'b1;
pika_color[3142] <= 1'b1;
pika_color[3179] <= 1'b1;
pika_color[3180] <= 1'b1;
pika_color[3195] <= 1'b1;
pika_color[3196] <= 1'b1;
pika_color[3197] <= 1'b1;
pika_color[3198] <= 1'b1;
pika_color[3229] <= 1'b1;
pika_color[3230] <= 1'b1;
pika_color[3231] <= 1'b1;
pika_color[3232] <= 1'b1;
pika_color[3233] <= 1'b1;
pika_color[3234] <= 1'b1;
pika_color[3235] <= 1'b1;
pika_color[3240] <= 1'b1;
pika_color[3241] <= 1'b1;
pika_color[3242] <= 1'b1;
pika_color[3243] <= 1'b1;
pika_color[3257] <= 1'b1;
pika_color[3258] <= 1'b1;
pika_color[3294] <= 1'b1;
pika_color[3310] <= 1'b1;
pika_color[3311] <= 1'b1;
pika_color[3312] <= 1'b1;
pika_color[3345] <= 1'b1;
pika_color[3346] <= 1'b1;
pika_color[3347] <= 1'b1;
pika_color[3348] <= 1'b1;
pika_color[3350] <= 1'b1;
pika_color[3357] <= 1'b1;
pika_color[3358] <= 1'b1;
pika_color[3359] <= 1'b1;
pika_color[3360] <= 1'b1;
pika_color[3373] <= 1'b1;
pika_color[3408] <= 1'b1;
pika_color[3409] <= 1'b1;
pika_color[3425] <= 1'b1;
pika_color[3426] <= 1'b1;
pika_color[3460] <= 1'b1;
pika_color[3461] <= 1'b1;
pika_color[3462] <= 1'b1;
pika_color[3463] <= 1'b1;
pika_color[3464] <= 1'b1;
pika_color[3465] <= 1'b1;
pika_color[3475] <= 1'b1;
pika_color[3476] <= 1'b1;
pika_color[3488] <= 1'b1;
pika_color[3489] <= 1'b1;
pika_color[3522] <= 1'b1;
pika_color[3523] <= 1'b1;
pika_color[3540] <= 1'b1;
pika_color[3576] <= 1'b1;
pika_color[3577] <= 1'b1;
pika_color[3578] <= 1'b1;
pika_color[3579] <= 1'b1;
pika_color[3580] <= 1'b1;
pika_color[3591] <= 1'b1;
pika_color[3604] <= 1'b1;
pika_color[3636] <= 1'b1;
pika_color[3637] <= 1'b1;
pika_color[3653] <= 1'b1;
pika_color[3654] <= 1'b1;
pika_color[3655] <= 1'b1;
pika_color[3691] <= 1'b1;
pika_color[3692] <= 1'b1;
pika_color[3693] <= 1'b1;
pika_color[3694] <= 1'b1;
pika_color[3695] <= 1'b1;
pika_color[3707] <= 1'b1;
pika_color[3708] <= 1'b1;
pika_color[3719] <= 1'b1;
pika_color[3720] <= 1'b1;
pika_color[3750] <= 1'b1;
pika_color[3751] <= 1'b1;
pika_color[3767] <= 1'b1;
pika_color[3768] <= 1'b1;
pika_color[3807] <= 1'b1;
pika_color[3808] <= 1'b1;
pika_color[3809] <= 1'b1;
pika_color[3810] <= 1'b1;
pika_color[3823] <= 1'b1;
pika_color[3824] <= 1'b1;
pika_color[3835] <= 1'b1;
pika_color[3865] <= 1'b1;
pika_color[3881] <= 1'b1;
pika_color[3882] <= 1'b1;
pika_color[3923] <= 1'b1;
pika_color[3924] <= 1'b1;
pika_color[3925] <= 1'b1;
pika_color[3939] <= 1'b1;
pika_color[3940] <= 1'b1;
pika_color[3941] <= 1'b1;
pika_color[3950] <= 1'b1;
pika_color[3951] <= 1'b1;
pika_color[3980] <= 1'b1;
pika_color[3996] <= 1'b1;
pika_color[4038] <= 1'b1;
pika_color[4039] <= 1'b1;
pika_color[4040] <= 1'b1;
pika_color[4056] <= 1'b1;
pika_color[4057] <= 1'b1;
pika_color[4067] <= 1'b1;
pika_color[4073] <= 1'b1;
pika_color[4074] <= 1'b1;
pika_color[4075] <= 1'b1;
pika_color[4076] <= 1'b1;
pika_color[4077] <= 1'b1;
pika_color[4078] <= 1'b1;
pika_color[4079] <= 1'b1;
pika_color[4080] <= 1'b1;
pika_color[4081] <= 1'b1;
pika_color[4082] <= 1'b1;
pika_color[4083] <= 1'b1;
pika_color[4084] <= 1'b1;
pika_color[4085] <= 1'b1;
pika_color[4086] <= 1'b1;
pika_color[4087] <= 1'b1;
pika_color[4088] <= 1'b1;
pika_color[4089] <= 1'b1;
pika_color[4094] <= 1'b1;
pika_color[4095] <= 1'b1;
pika_color[4110] <= 1'b1;
pika_color[4111] <= 1'b1;
pika_color[4154] <= 1'b1;
pika_color[4155] <= 1'b1;
pika_color[4172] <= 1'b1;
pika_color[4173] <= 1'b1;
pika_color[4182] <= 1'b1;
pika_color[4185] <= 1'b1;
pika_color[4186] <= 1'b1;
pika_color[4187] <= 1'b1;
pika_color[4188] <= 1'b1;
pika_color[4204] <= 1'b1;
pika_color[4205] <= 1'b1;
pika_color[4206] <= 1'b1;
pika_color[4208] <= 1'b1;
pika_color[4209] <= 1'b1;
pika_color[4223] <= 1'b1;
pika_color[4224] <= 1'b1;
pika_color[4225] <= 1'b1;
pika_color[4270] <= 1'b1;
pika_color[4271] <= 1'b1;
pika_color[4288] <= 1'b1;
pika_color[4289] <= 1'b1;
pika_color[4297] <= 1'b1;
pika_color[4298] <= 1'b1;
pika_color[4299] <= 1'b1;
pika_color[4300] <= 1'b1;
pika_color[4322] <= 1'b1;
pika_color[4323] <= 1'b1;
pika_color[4337] <= 1'b1;
pika_color[4338] <= 1'b1;
pika_color[4386] <= 1'b1;
pika_color[4387] <= 1'b1;
pika_color[4404] <= 1'b1;
pika_color[4405] <= 1'b1;
pika_color[4412] <= 1'b1;
pika_color[4413] <= 1'b1;
pika_color[4451] <= 1'b1;
pika_color[4452] <= 1'b1;
pika_color[4502] <= 1'b1;
pika_color[4503] <= 1'b1;
pika_color[4520] <= 1'b1;
pika_color[4521] <= 1'b1;
pika_color[4526] <= 1'b1;
pika_color[4527] <= 1'b1;
pika_color[4564] <= 1'b1;
pika_color[4565] <= 1'b1;
pika_color[4566] <= 1'b1;
pika_color[4618] <= 1'b1;
pika_color[4619] <= 1'b1;
pika_color[4636] <= 1'b1;
pika_color[4637] <= 1'b1;
pika_color[4639] <= 1'b1;
pika_color[4640] <= 1'b1;
pika_color[4677] <= 1'b1;
pika_color[4678] <= 1'b1;
pika_color[4679] <= 1'b1;
pika_color[4734] <= 1'b1;
pika_color[4752] <= 1'b1;
pika_color[4753] <= 1'b1;
pika_color[4754] <= 1'b1;
pika_color[4791] <= 1'b1;
pika_color[4792] <= 1'b1;
pika_color[4850] <= 1'b1;
pika_color[4867] <= 1'b1;
pika_color[4868] <= 1'b1;
pika_color[4869] <= 1'b1;
pika_color[4905] <= 1'b1;
pika_color[4906] <= 1'b1;
pika_color[4965] <= 1'b1;
pika_color[4966] <= 1'b1;
pika_color[4984] <= 1'b1;
pika_color[5021] <= 1'b1;
pika_color[5081] <= 1'b1;
pika_color[5082] <= 1'b1;
pika_color[5099] <= 1'b1;
pika_color[5136] <= 1'b1;
pika_color[5137] <= 1'b1;
pika_color[5197] <= 1'b1;
pika_color[5198] <= 1'b1;
pika_color[5252] <= 1'b1;
pika_color[5313] <= 1'b1;
pika_color[5314] <= 1'b1;
pika_color[5315] <= 1'b1;
pika_color[5367] <= 1'b1;
pika_color[5368] <= 1'b1;
pika_color[5430] <= 1'b1;
pika_color[5431] <= 1'b1;
pika_color[5483] <= 1'b1;
pika_color[5546] <= 1'b1;
pika_color[5547] <= 1'b1;
pika_color[5598] <= 1'b1;
pika_color[5599] <= 1'b1;
pika_color[5662] <= 1'b1;
pika_color[5663] <= 1'b1;
pika_color[5715] <= 1'b1;
pika_color[5779] <= 1'b1;
pika_color[5780] <= 1'b1;
pika_color[5781] <= 1'b1;
pika_color[5830] <= 1'b1;
pika_color[5831] <= 1'b1;
pika_color[5896] <= 1'b1;
pika_color[5897] <= 1'b1;
pika_color[5946] <= 1'b1;
pika_color[6012] <= 1'b1;
pika_color[6013] <= 1'b1;
pika_color[6061] <= 1'b1;
pika_color[6127] <= 1'b1;
pika_color[6176] <= 1'b1;
pika_color[6177] <= 1'b1;
pika_color[6242] <= 1'b1;
pika_color[6292] <= 1'b1;
pika_color[6357] <= 1'b1;
pika_color[6407] <= 1'b1;
pika_color[6472] <= 1'b1;
pika_color[6522] <= 1'b1;
pika_color[6587] <= 1'b1;
pika_color[6622] <= 1'b1;
pika_color[6623] <= 1'b1;
pika_color[6624] <= 1'b1;
pika_color[6625] <= 1'b1;
pika_color[6637] <= 1'b1;
pika_color[6638] <= 1'b1;
pika_color[6702] <= 1'b1;
pika_color[6735] <= 1'b1;
pika_color[6736] <= 1'b1;
pika_color[6737] <= 1'b1;
pika_color[6738] <= 1'b1;
pika_color[6739] <= 1'b1;
pika_color[6753] <= 1'b1;
pika_color[6817] <= 1'b1;
pika_color[6850] <= 1'b1;
pika_color[6851] <= 1'b1;
pika_color[6864] <= 1'b1;
pika_color[6865] <= 1'b1;
pika_color[6866] <= 1'b1;
pika_color[6867] <= 1'b1;
pika_color[6868] <= 1'b1;
pika_color[6932] <= 1'b1;
pika_color[6979] <= 1'b1;
pika_color[6983] <= 1'b1;
pika_color[6984] <= 1'b1;
pika_color[6985] <= 1'b1;
pika_color[7047] <= 1'b1;
pika_color[7093] <= 1'b1;
pika_color[7101] <= 1'b1;
pika_color[7102] <= 1'b1;
pika_color[7162] <= 1'b1;
pika_color[7208] <= 1'b1;
pika_color[7217] <= 1'b1;
pika_color[7277] <= 1'b1;
pika_color[7287] <= 1'b1;
pika_color[7288] <= 1'b1;
pika_color[7289] <= 1'b1;
pika_color[7290] <= 1'b1;
pika_color[7291] <= 1'b1;
pika_color[7292] <= 1'b1;
pika_color[7293] <= 1'b1;
pika_color[7323] <= 1'b1;
pika_color[7332] <= 1'b1;
pika_color[7333] <= 1'b1;
pika_color[7392] <= 1'b1;
pika_color[7401] <= 1'b1;
pika_color[7402] <= 1'b1;
pika_color[7403] <= 1'b1;
pika_color[7404] <= 1'b1;
pika_color[7405] <= 1'b1;
pika_color[7406] <= 1'b1;
pika_color[7407] <= 1'b1;
pika_color[7408] <= 1'b1;
pika_color[7438] <= 1'b1;
pika_color[7448] <= 1'b1;
pika_color[7449] <= 1'b1;
pika_color[7507] <= 1'b1;
pika_color[7531] <= 1'b1;
pika_color[7532] <= 1'b1;
pika_color[7533] <= 1'b1;
pika_color[7534] <= 1'b1;
pika_color[7535] <= 1'b1;
pika_color[7553] <= 1'b1;
pika_color[7554] <= 1'b1;
pika_color[7564] <= 1'b1;
pika_color[7622] <= 1'b1;
pika_color[7645] <= 1'b1;
pika_color[7646] <= 1'b1;
pika_color[7647] <= 1'b1;
pika_color[7648] <= 1'b1;
pika_color[7649] <= 1'b1;
pika_color[7669] <= 1'b1;
pika_color[7679] <= 1'b1;
pika_color[7737] <= 1'b1;
pika_color[7761] <= 1'b1;
pika_color[7762] <= 1'b1;
pika_color[7763] <= 1'b1;
pika_color[7784] <= 1'b1;
pika_color[7794] <= 1'b1;
pika_color[7795] <= 1'b1;
pika_color[7852] <= 1'b1;
pika_color[7899] <= 1'b1;
pika_color[7910] <= 1'b1;
pika_color[7967] <= 1'b1;
pika_color[8013] <= 1'b1;
pika_color[8014] <= 1'b1;
pika_color[8025] <= 1'b1;
pika_color[8082] <= 1'b1;
pika_color[8083] <= 1'b1;
pika_color[8128] <= 1'b1;
pika_color[8140] <= 1'b1;
pika_color[8198] <= 1'b1;
pika_color[8220] <= 1'b1;
pika_color[8221] <= 1'b1;
pika_color[8222] <= 1'b1;
pika_color[8223] <= 1'b1;
pika_color[8224] <= 1'b1;
pika_color[8225] <= 1'b1;
pika_color[8226] <= 1'b1;
pika_color[8227] <= 1'b1;
pika_color[8228] <= 1'b1;
pika_color[8229] <= 1'b1;
pika_color[8243] <= 1'b1;
pika_color[8255] <= 1'b1;
pika_color[8313] <= 1'b1;
pika_color[8334] <= 1'b1;
pika_color[8335] <= 1'b1;
pika_color[8344] <= 1'b1;
pika_color[8357] <= 1'b1;
pika_color[8358] <= 1'b1;
pika_color[8370] <= 1'b1;
pika_color[8428] <= 1'b1;
pika_color[8447] <= 1'b1;
pika_color[8448] <= 1'b1;
pika_color[8452] <= 1'b1;
pika_color[8453] <= 1'b1;
pika_color[8454] <= 1'b1;
pika_color[8455] <= 1'b1;
pika_color[8456] <= 1'b1;
pika_color[8457] <= 1'b1;
pika_color[8458] <= 1'b1;
pika_color[8459] <= 1'b1;
pika_color[8472] <= 1'b1;
pika_color[8485] <= 1'b1;
pika_color[8543] <= 1'b1;
pika_color[8544] <= 1'b1;
pika_color[8562] <= 1'b1;
pika_color[8563] <= 1'b1;
pika_color[8565] <= 1'b1;
pika_color[8566] <= 1'b1;
pika_color[8567] <= 1'b1;
pika_color[8573] <= 1'b1;
pika_color[8586] <= 1'b1;
pika_color[8587] <= 1'b1;
pika_color[8600] <= 1'b1;
pika_color[8659] <= 1'b1;
pika_color[8678] <= 1'b1;
pika_color[8679] <= 1'b1;
pika_color[8680] <= 1'b1;
pika_color[8687] <= 1'b1;
pika_color[8688] <= 1'b1;
pika_color[8701] <= 1'b1;
pika_color[8715] <= 1'b1;
pika_color[8774] <= 1'b1;
pika_color[8775] <= 1'b1;
pika_color[8794] <= 1'b1;
pika_color[8795] <= 1'b1;
pika_color[8801] <= 1'b1;
pika_color[8802] <= 1'b1;
pika_color[8815] <= 1'b1;
pika_color[8816] <= 1'b1;
pika_color[8830] <= 1'b1;
pika_color[8890] <= 1'b1;
pika_color[8910] <= 1'b1;
pika_color[8911] <= 1'b1;
pika_color[8912] <= 1'b1;
pika_color[8913] <= 1'b1;
pika_color[8914] <= 1'b1;
pika_color[8915] <= 1'b1;
pika_color[8916] <= 1'b1;
pika_color[8930] <= 1'b1;
pika_color[8945] <= 1'b1;
pika_color[9005] <= 1'b1;
pika_color[9006] <= 1'b1;
pika_color[9044] <= 1'b1;
pika_color[9045] <= 1'b1;
pika_color[9060] <= 1'b1;
pika_color[9121] <= 1'b1;
pika_color[9122] <= 1'b1;
pika_color[9159] <= 1'b1;
pika_color[9175] <= 1'b1;
pika_color[9236] <= 1'b1;
pika_color[9237] <= 1'b1;
pika_color[9238] <= 1'b1;
pika_color[9274] <= 1'b1;
pika_color[9290] <= 1'b1;
pika_color[9350] <= 1'b1;
pika_color[9351] <= 1'b1;
pika_color[9353] <= 1'b1;
pika_color[9354] <= 1'b1;
pika_color[9388] <= 1'b1;
pika_color[9405] <= 1'b1;
pika_color[9465] <= 1'b1;
pika_color[9469] <= 1'b1;
pika_color[9470] <= 1'b1;
pika_color[9471] <= 1'b1;
pika_color[9502] <= 1'b1;
pika_color[9503] <= 1'b1;
pika_color[9520] <= 1'b1;
pika_color[9579] <= 1'b1;
pika_color[9580] <= 1'b1;
pika_color[9586] <= 1'b1;
pika_color[9587] <= 1'b1;
pika_color[9617] <= 1'b1;
pika_color[9635] <= 1'b1;
pika_color[9693] <= 1'b1;
pika_color[9694] <= 1'b1;
pika_color[9703] <= 1'b1;
pika_color[9704] <= 1'b1;
pika_color[9705] <= 1'b1;
pika_color[9732] <= 1'b1;
pika_color[9750] <= 1'b1;
pika_color[9808] <= 1'b1;
pika_color[9846] <= 1'b1;
pika_color[9847] <= 1'b1;
pika_color[9865] <= 1'b1;
pika_color[9922] <= 1'b1;
pika_color[9923] <= 1'b1;
pika_color[9936] <= 1'b1;
pika_color[9937] <= 1'b1;
pika_color[9960] <= 1'b1;
pika_color[9961] <= 1'b1;
pika_color[9980] <= 1'b1;
pika_color[10037] <= 1'b1;
pika_color[10050] <= 1'b1;
pika_color[10051] <= 1'b1;
pika_color[10095] <= 1'b1;
pika_color[10152] <= 1'b1;
pika_color[10165] <= 1'b1;
pika_color[10210] <= 1'b1;
pika_color[10267] <= 1'b1;
pika_color[10280] <= 1'b1;
pika_color[10325] <= 1'b1;
pika_color[10382] <= 1'b1;
pika_color[10395] <= 1'b1;
pika_color[10396] <= 1'b1;
pika_color[10440] <= 1'b1;
pika_color[10497] <= 1'b1;
pika_color[10511] <= 1'b1;
pika_color[10512] <= 1'b1;
pika_color[10555] <= 1'b1;
pika_color[10612] <= 1'b1;
pika_color[10627] <= 1'b1;
pika_color[10670] <= 1'b1;
pika_color[10727] <= 1'b1;
pika_color[10742] <= 1'b1;
pika_color[10743] <= 1'b1;
pika_color[10785] <= 1'b1;
pika_color[10842] <= 1'b1;
pika_color[10858] <= 1'b1;
pika_color[10900] <= 1'b1;
pika_color[10957] <= 1'b1;
pika_color[10958] <= 1'b1;
pika_color[10973] <= 1'b1;
pika_color[11015] <= 1'b1;
pika_color[11073] <= 1'b1;
pika_color[11088] <= 1'b1;
pika_color[11130] <= 1'b1;
pika_color[11188] <= 1'b1;
pika_color[11189] <= 1'b1;
pika_color[11202] <= 1'b1;
pika_color[11203] <= 1'b1;
pika_color[11245] <= 1'b1;
pika_color[11304] <= 1'b1;
pika_color[11317] <= 1'b1;
pika_color[11360] <= 1'b1;
pika_color[11419] <= 1'b1;
pika_color[11420] <= 1'b1;
pika_color[11431] <= 1'b1;
pika_color[11432] <= 1'b1;
pika_color[11475] <= 1'b1;
pika_color[11535] <= 1'b1;
pika_color[11545] <= 1'b1;
pika_color[11546] <= 1'b1;
pika_color[11590] <= 1'b1;
pika_color[11650] <= 1'b1;
pika_color[11651] <= 1'b1;
pika_color[11660] <= 1'b1;
pika_color[11705] <= 1'b1;
pika_color[11706] <= 1'b1;
pika_color[11765] <= 1'b1;
pika_color[11766] <= 1'b1;
pika_color[11767] <= 1'b1;
pika_color[11768] <= 1'b1;
pika_color[11769] <= 1'b1;
pika_color[11773] <= 1'b1;
pika_color[11774] <= 1'b1;
pika_color[11775] <= 1'b1;
pika_color[11821] <= 1'b1;
pika_color[11880] <= 1'b1;
pika_color[11884] <= 1'b1;
pika_color[11885] <= 1'b1;
pika_color[11886] <= 1'b1;
pika_color[11887] <= 1'b1;
pika_color[11888] <= 1'b1;
pika_color[11936] <= 1'b1;
pika_color[11995] <= 1'b1;
pika_color[12051] <= 1'b1;
pika_color[12110] <= 1'b1;
pika_color[12166] <= 1'b1;
pika_color[12225] <= 1'b1;
pika_color[12281] <= 1'b1;
pika_color[12282] <= 1'b1;
pika_color[12340] <= 1'b1;
pika_color[12397] <= 1'b1;
pika_color[12455] <= 1'b1;
pika_color[12512] <= 1'b1;
pika_color[12570] <= 1'b1;
pika_color[12627] <= 1'b1;
pika_color[12685] <= 1'b1;
pika_color[12742] <= 1'b1;
pika_color[12800] <= 1'b1;
pika_color[12857] <= 1'b1;
pika_color[12915] <= 1'b1;
pika_color[12972] <= 1'b1;
pika_color[13030] <= 1'b1;
pika_color[13087] <= 1'b1;
pika_color[13145] <= 1'b1;
pika_color[13202] <= 1'b1;
pika_color[13260] <= 1'b1;
pika_color[13317] <= 1'b1;
pika_color[13375] <= 1'b1;
pika_color[13376] <= 1'b1;
pika_color[13432] <= 1'b1;
pika_color[13491] <= 1'b1;
pika_color[13547] <= 1'b1;
pika_color[13606] <= 1'b1;
pika_color[13662] <= 1'b1;
pika_color[13721] <= 1'b1;
pika_color[13722] <= 1'b1;
pika_color[13777] <= 1'b1;
pika_color[13837] <= 1'b1;
pika_color[13892] <= 1'b1;
pika_color[13952] <= 1'b1;
pika_color[14007] <= 1'b1;
pika_color[14067] <= 1'b1;
pika_color[14122] <= 1'b1;
pika_color[14182] <= 1'b1;
pika_color[14183] <= 1'b1;
pika_color[14237] <= 1'b1;
pika_color[14298] <= 1'b1;
pika_color[14352] <= 1'b1;
pika_color[14413] <= 1'b1;
pika_color[14414] <= 1'b1;
pika_color[14466] <= 1'b1;
pika_color[14467] <= 1'b1;
pika_color[14529] <= 1'b1;
pika_color[14581] <= 1'b1;
pika_color[14644] <= 1'b1;
pika_color[14645] <= 1'b1;
pika_color[14695] <= 1'b1;
pika_color[14696] <= 1'b1;
pika_color[14760] <= 1'b1;
pika_color[14810] <= 1'b1;
pika_color[14876] <= 1'b1;
pika_color[14925] <= 1'b1;
pika_color[14991] <= 1'b1;
pika_color[14992] <= 1'b1;
pika_color[15039] <= 1'b1;
pika_color[15040] <= 1'b1;
pika_color[15107] <= 1'b1;
pika_color[15108] <= 1'b1;
pika_color[15154] <= 1'b1;
pika_color[15223] <= 1'b1;
pika_color[15224] <= 1'b1;
pika_color[15267] <= 1'b1;
pika_color[15268] <= 1'b1;
pika_color[15269] <= 1'b1;
pika_color[15339] <= 1'b1;
pika_color[15340] <= 1'b1;
pika_color[15341] <= 1'b1;
pika_color[15353] <= 1'b1;
pika_color[15354] <= 1'b1;
pika_color[15355] <= 1'b1;
pika_color[15356] <= 1'b1;
pika_color[15357] <= 1'b1;
pika_color[15358] <= 1'b1;
pika_color[15359] <= 1'b1;
pika_color[15382] <= 1'b1;
pika_color[15456] <= 1'b1;
pika_color[15457] <= 1'b1;
pika_color[15458] <= 1'b1;
pika_color[15468] <= 1'b1;
pika_color[15474] <= 1'b1;
pika_color[15475] <= 1'b1;
pika_color[15476] <= 1'b1;
pika_color[15477] <= 1'b1;
pika_color[15478] <= 1'b1;
pika_color[15496] <= 1'b1;
pika_color[15497] <= 1'b1;
pika_color[15573] <= 1'b1;
pika_color[15574] <= 1'b1;
pika_color[15583] <= 1'b1;
pika_color[15593] <= 1'b1;
pika_color[15594] <= 1'b1;
pika_color[15595] <= 1'b1;
pika_color[15596] <= 1'b1;
pika_color[15597] <= 1'b1;
pika_color[15610] <= 1'b1;
pika_color[15611] <= 1'b1;
pika_color[15689] <= 1'b1;
pika_color[15697] <= 1'b1;
pika_color[15698] <= 1'b1;
pika_color[15712] <= 1'b1;
pika_color[15713] <= 1'b1;
pika_color[15722] <= 1'b1;
pika_color[15723] <= 1'b1;
pika_color[15724] <= 1'b1;
pika_color[15725] <= 1'b1;
pika_color[15804] <= 1'b1;
pika_color[15805] <= 1'b1;
pika_color[15812] <= 1'b1;
pika_color[15828] <= 1'b1;
pika_color[15836] <= 1'b1;
pika_color[15837] <= 1'b1;
pika_color[15921] <= 1'b1;
pika_color[15922] <= 1'b1;
pika_color[15923] <= 1'b1;
pika_color[15924] <= 1'b1;
pika_color[15925] <= 1'b1;
pika_color[15926] <= 1'b1;
pika_color[15942] <= 1'b1;
pika_color[15943] <= 1'b1;
pika_color[15951] <= 1'b1;
pika_color[16057] <= 1'b1;
pika_color[16066] <= 1'b1;
pika_color[16172] <= 1'b1;
pika_color[16181] <= 1'b1;
pika_color[16287] <= 1'b1;
pika_color[16288] <= 1'b1;
pika_color[16289] <= 1'b1;
pika_color[16290] <= 1'b1;
pika_color[16291] <= 1'b1;
pika_color[16292] <= 1'b1;
pika_color[16293] <= 1'b1;
pika_color[16294] <= 1'b1;
pika_color[16295] <= 1'b1;
pika_color[16296] <= 1'b1;


		end
		move50, move51, move52, move53, move54, move55, move56, move57, move58, move59:
		begin
		
pika_color[890] <= 1'b1;
pika_color[891] <= 1'b1;
pika_color[892] <= 1'b1;
pika_color[893] <= 1'b1;
pika_color[894] <= 1'b1;
pika_color[895] <= 1'b1;
pika_color[896] <= 1'b1;
pika_color[897] <= 1'b1;
pika_color[1002] <= 1'b1;
pika_color[1003] <= 1'b1;
pika_color[1004] <= 1'b1;
pika_color[1005] <= 1'b1;
pika_color[1006] <= 1'b1;
pika_color[1007] <= 1'b1;
pika_color[1008] <= 1'b1;
pika_color[1009] <= 1'b1;
pika_color[1010] <= 1'b1;
pika_color[1011] <= 1'b1;
pika_color[1012] <= 1'b1;
pika_color[1116] <= 1'b1;
pika_color[1117] <= 1'b1;
pika_color[1120] <= 1'b1;
pika_color[1121] <= 1'b1;
pika_color[1122] <= 1'b1;
pika_color[1123] <= 1'b1;
pika_color[1124] <= 1'b1;
pika_color[1125] <= 1'b1;
pika_color[1126] <= 1'b1;
pika_color[1127] <= 1'b1;
pika_color[1229] <= 1'b1;
pika_color[1230] <= 1'b1;
pika_color[1235] <= 1'b1;
pika_color[1236] <= 1'b1;
pika_color[1237] <= 1'b1;
pika_color[1238] <= 1'b1;
pika_color[1239] <= 1'b1;
pika_color[1240] <= 1'b1;
pika_color[1241] <= 1'b1;
pika_color[1242] <= 1'b1;
pika_color[1342] <= 1'b1;
pika_color[1343] <= 1'b1;
pika_color[1344] <= 1'b1;
pika_color[1350] <= 1'b1;
pika_color[1351] <= 1'b1;
pika_color[1352] <= 1'b1;
pika_color[1353] <= 1'b1;
pika_color[1354] <= 1'b1;
pika_color[1355] <= 1'b1;
pika_color[1356] <= 1'b1;
pika_color[1357] <= 1'b1;
pika_color[1389] <= 1'b1;
pika_color[1390] <= 1'b1;
pika_color[1391] <= 1'b1;
pika_color[1392] <= 1'b1;
pika_color[1393] <= 1'b1;
pika_color[1394] <= 1'b1;
pika_color[1456] <= 1'b1;
pika_color[1457] <= 1'b1;
pika_color[1465] <= 1'b1;
pika_color[1466] <= 1'b1;
pika_color[1467] <= 1'b1;
pika_color[1468] <= 1'b1;
pika_color[1469] <= 1'b1;
pika_color[1470] <= 1'b1;
pika_color[1471] <= 1'b1;
pika_color[1504] <= 1'b1;
pika_color[1505] <= 1'b1;
pika_color[1506] <= 1'b1;
pika_color[1507] <= 1'b1;
pika_color[1508] <= 1'b1;
pika_color[1509] <= 1'b1;
pika_color[1510] <= 1'b1;
pika_color[1511] <= 1'b1;
pika_color[1570] <= 1'b1;
pika_color[1571] <= 1'b1;
pika_color[1580] <= 1'b1;
pika_color[1581] <= 1'b1;
pika_color[1582] <= 1'b1;
pika_color[1583] <= 1'b1;
pika_color[1584] <= 1'b1;
pika_color[1585] <= 1'b1;
pika_color[1586] <= 1'b1;
pika_color[1619] <= 1'b1;
pika_color[1620] <= 1'b1;
pika_color[1621] <= 1'b1;
pika_color[1622] <= 1'b1;
pika_color[1623] <= 1'b1;
pika_color[1624] <= 1'b1;
pika_color[1625] <= 1'b1;
pika_color[1626] <= 1'b1;
pika_color[1627] <= 1'b1;
pika_color[1628] <= 1'b1;
pika_color[1684] <= 1'b1;
pika_color[1685] <= 1'b1;
pika_color[1695] <= 1'b1;
pika_color[1696] <= 1'b1;
pika_color[1697] <= 1'b1;
pika_color[1698] <= 1'b1;
pika_color[1699] <= 1'b1;
pika_color[1700] <= 1'b1;
pika_color[1734] <= 1'b1;
pika_color[1735] <= 1'b1;
pika_color[1736] <= 1'b1;
pika_color[1737] <= 1'b1;
pika_color[1738] <= 1'b1;
pika_color[1739] <= 1'b1;
pika_color[1740] <= 1'b1;
pika_color[1743] <= 1'b1;
pika_color[1744] <= 1'b1;
pika_color[1745] <= 1'b1;
pika_color[1798] <= 1'b1;
pika_color[1799] <= 1'b1;
pika_color[1810] <= 1'b1;
pika_color[1811] <= 1'b1;
pika_color[1812] <= 1'b1;
pika_color[1813] <= 1'b1;
pika_color[1814] <= 1'b1;
pika_color[1815] <= 1'b1;
pika_color[1849] <= 1'b1;
pika_color[1850] <= 1'b1;
pika_color[1851] <= 1'b1;
pika_color[1852] <= 1'b1;
pika_color[1853] <= 1'b1;
pika_color[1854] <= 1'b1;
pika_color[1855] <= 1'b1;
pika_color[1860] <= 1'b1;
pika_color[1861] <= 1'b1;
pika_color[1862] <= 1'b1;
pika_color[1912] <= 1'b1;
pika_color[1913] <= 1'b1;
pika_color[1925] <= 1'b1;
pika_color[1926] <= 1'b1;
pika_color[1927] <= 1'b1;
pika_color[1928] <= 1'b1;
pika_color[1929] <= 1'b1;
pika_color[1965] <= 1'b1;
pika_color[1966] <= 1'b1;
pika_color[1967] <= 1'b1;
pika_color[1968] <= 1'b1;
pika_color[1969] <= 1'b1;
pika_color[1970] <= 1'b1;
pika_color[1976] <= 1'b1;
pika_color[1977] <= 1'b1;
pika_color[1978] <= 1'b1;
pika_color[2026] <= 1'b1;
pika_color[2027] <= 1'b1;
pika_color[2040] <= 1'b1;
pika_color[2041] <= 1'b1;
pika_color[2042] <= 1'b1;
pika_color[2043] <= 1'b1;
pika_color[2080] <= 1'b1;
pika_color[2081] <= 1'b1;
pika_color[2082] <= 1'b1;
pika_color[2083] <= 1'b1;
pika_color[2084] <= 1'b1;
pika_color[2085] <= 1'b1;
pika_color[2093] <= 1'b1;
pika_color[2094] <= 1'b1;
pika_color[2141] <= 1'b1;
pika_color[2155] <= 1'b1;
pika_color[2156] <= 1'b1;
pika_color[2157] <= 1'b1;
pika_color[2195] <= 1'b1;
pika_color[2196] <= 1'b1;
pika_color[2197] <= 1'b1;
pika_color[2198] <= 1'b1;
pika_color[2199] <= 1'b1;
pika_color[2200] <= 1'b1;
pika_color[2209] <= 1'b1;
pika_color[2210] <= 1'b1;
pika_color[2255] <= 1'b1;
pika_color[2270] <= 1'b1;
pika_color[2271] <= 1'b1;
pika_color[2272] <= 1'b1;
pika_color[2311] <= 1'b1;
pika_color[2312] <= 1'b1;
pika_color[2313] <= 1'b1;
pika_color[2314] <= 1'b1;
pika_color[2315] <= 1'b1;
pika_color[2325] <= 1'b1;
pika_color[2369] <= 1'b1;
pika_color[2370] <= 1'b1;
pika_color[2385] <= 1'b1;
pika_color[2386] <= 1'b1;
pika_color[2426] <= 1'b1;
pika_color[2427] <= 1'b1;
pika_color[2428] <= 1'b1;
pika_color[2429] <= 1'b1;
pika_color[2430] <= 1'b1;
pika_color[2440] <= 1'b1;
pika_color[2441] <= 1'b1;
pika_color[2483] <= 1'b1;
pika_color[2484] <= 1'b1;
pika_color[2500] <= 1'b1;
pika_color[2542] <= 1'b1;
pika_color[2543] <= 1'b1;
pika_color[2544] <= 1'b1;
pika_color[2545] <= 1'b1;
pika_color[2556] <= 1'b1;
pika_color[2557] <= 1'b1;
pika_color[2558] <= 1'b1;
pika_color[2598] <= 1'b1;
pika_color[2615] <= 1'b1;
pika_color[2657] <= 1'b1;
pika_color[2658] <= 1'b1;
pika_color[2659] <= 1'b1;
pika_color[2660] <= 1'b1;
pika_color[2673] <= 1'b1;
pika_color[2674] <= 1'b1;
pika_color[2712] <= 1'b1;
pika_color[2713] <= 1'b1;
pika_color[2729] <= 1'b1;
pika_color[2730] <= 1'b1;
pika_color[2773] <= 1'b1;
pika_color[2774] <= 1'b1;
pika_color[2775] <= 1'b1;
pika_color[2789] <= 1'b1;
pika_color[2790] <= 1'b1;
pika_color[2826] <= 1'b1;
pika_color[2827] <= 1'b1;
pika_color[2843] <= 1'b1;
pika_color[2844] <= 1'b1;
pika_color[2888] <= 1'b1;
pika_color[2889] <= 1'b1;
pika_color[2890] <= 1'b1;
pika_color[2905] <= 1'b1;
pika_color[2906] <= 1'b1;
pika_color[2941] <= 1'b1;
pika_color[2958] <= 1'b1;
pika_color[3004] <= 1'b1;
pika_color[3005] <= 1'b1;
pika_color[3020] <= 1'b1;
pika_color[3021] <= 1'b1;
pika_color[3055] <= 1'b1;
pika_color[3056] <= 1'b1;
pika_color[3072] <= 1'b1;
pika_color[3073] <= 1'b1;
pika_color[3120] <= 1'b1;
pika_color[3136] <= 1'b1;
pika_color[3137] <= 1'b1;
pika_color[3170] <= 1'b1;
pika_color[3186] <= 1'b1;
pika_color[3187] <= 1'b1;
pika_color[3235] <= 1'b1;
pika_color[3236] <= 1'b1;
pika_color[3252] <= 1'b1;
pika_color[3267] <= 1'b1;
pika_color[3268] <= 1'b1;
pika_color[3269] <= 1'b1;
pika_color[3270] <= 1'b1;
pika_color[3271] <= 1'b1;
pika_color[3272] <= 1'b1;
pika_color[3273] <= 1'b1;
pika_color[3274] <= 1'b1;
pika_color[3275] <= 1'b1;
pika_color[3276] <= 1'b1;
pika_color[3277] <= 1'b1;
pika_color[3278] <= 1'b1;
pika_color[3279] <= 1'b1;
pika_color[3284] <= 1'b1;
pika_color[3300] <= 1'b1;
pika_color[3301] <= 1'b1;
pika_color[3351] <= 1'b1;
pika_color[3352] <= 1'b1;
pika_color[3368] <= 1'b1;
pika_color[3378] <= 1'b1;
pika_color[3379] <= 1'b1;
pika_color[3380] <= 1'b1;
pika_color[3381] <= 1'b1;
pika_color[3382] <= 1'b1;
pika_color[3394] <= 1'b1;
pika_color[3395] <= 1'b1;
pika_color[3396] <= 1'b1;
pika_color[3398] <= 1'b1;
pika_color[3413] <= 1'b1;
pika_color[3414] <= 1'b1;
pika_color[3415] <= 1'b1;
pika_color[3467] <= 1'b1;
pika_color[3483] <= 1'b1;
pika_color[3484] <= 1'b1;
pika_color[3491] <= 1'b1;
pika_color[3492] <= 1'b1;
pika_color[3493] <= 1'b1;
pika_color[3511] <= 1'b1;
pika_color[3512] <= 1'b1;
pika_color[3513] <= 1'b1;
pika_color[3527] <= 1'b1;
pika_color[3528] <= 1'b1;
pika_color[3582] <= 1'b1;
pika_color[3583] <= 1'b1;
pika_color[3599] <= 1'b1;
pika_color[3604] <= 1'b1;
pika_color[3605] <= 1'b1;
pika_color[3606] <= 1'b1;
pika_color[3641] <= 1'b1;
pika_color[3642] <= 1'b1;
pika_color[3698] <= 1'b1;
pika_color[3714] <= 1'b1;
pika_color[3715] <= 1'b1;
pika_color[3716] <= 1'b1;
pika_color[3717] <= 1'b1;
pika_color[3718] <= 1'b1;
pika_color[3719] <= 1'b1;
pika_color[3755] <= 1'b1;
pika_color[3756] <= 1'b1;
pika_color[3813] <= 1'b1;
pika_color[3814] <= 1'b1;
pika_color[3830] <= 1'b1;
pika_color[3831] <= 1'b1;
pika_color[3869] <= 1'b1;
pika_color[3870] <= 1'b1;
pika_color[3928] <= 1'b1;
pika_color[3929] <= 1'b1;
pika_color[3930] <= 1'b1;
pika_color[3946] <= 1'b1;
pika_color[3947] <= 1'b1;
pika_color[3983] <= 1'b1;
pika_color[3984] <= 1'b1;
pika_color[4044] <= 1'b1;
pika_color[4045] <= 1'b1;
pika_color[4046] <= 1'b1;
pika_color[4062] <= 1'b1;
pika_color[4097] <= 1'b1;
pika_color[4098] <= 1'b1;
pika_color[4159] <= 1'b1;
pika_color[4161] <= 1'b1;
pika_color[4162] <= 1'b1;
pika_color[4177] <= 1'b1;
pika_color[4178] <= 1'b1;
pika_color[4212] <= 1'b1;
pika_color[4213] <= 1'b1;
pika_color[4274] <= 1'b1;
pika_color[4275] <= 1'b1;
pika_color[4277] <= 1'b1;
pika_color[4278] <= 1'b1;
pika_color[4293] <= 1'b1;
pika_color[4328] <= 1'b1;
pika_color[4329] <= 1'b1;
pika_color[4390] <= 1'b1;
pika_color[4393] <= 1'b1;
pika_color[4394] <= 1'b1;
pika_color[4444] <= 1'b1;
pika_color[4505] <= 1'b1;
pika_color[4506] <= 1'b1;
pika_color[4509] <= 1'b1;
pika_color[4510] <= 1'b1;
pika_color[4559] <= 1'b1;
pika_color[4621] <= 1'b1;
pika_color[4625] <= 1'b1;
pika_color[4626] <= 1'b1;
pika_color[4674] <= 1'b1;
pika_color[4675] <= 1'b1;
pika_color[4736] <= 1'b1;
pika_color[4737] <= 1'b1;
pika_color[4741] <= 1'b1;
pika_color[4790] <= 1'b1;
pika_color[4852] <= 1'b1;
pika_color[4857] <= 1'b1;
pika_color[4906] <= 1'b1;
pika_color[4967] <= 1'b1;
pika_color[4972] <= 1'b1;
pika_color[4973] <= 1'b1;
pika_color[4974] <= 1'b1;
pika_color[5021] <= 1'b1;
pika_color[5022] <= 1'b1;
pika_color[5082] <= 1'b1;
pika_color[5083] <= 1'b1;
pika_color[5088] <= 1'b1;
pika_color[5089] <= 1'b1;
pika_color[5090] <= 1'b1;
pika_color[5137] <= 1'b1;
pika_color[5198] <= 1'b1;
pika_color[5203] <= 1'b1;
pika_color[5205] <= 1'b1;
pika_color[5206] <= 1'b1;
pika_color[5252] <= 1'b1;
pika_color[5253] <= 1'b1;
pika_color[5313] <= 1'b1;
pika_color[5314] <= 1'b1;
pika_color[5318] <= 1'b1;
pika_color[5321] <= 1'b1;
pika_color[5368] <= 1'b1;
pika_color[5429] <= 1'b1;
pika_color[5433] <= 1'b1;
pika_color[5483] <= 1'b1;
pika_color[5544] <= 1'b1;
pika_color[5545] <= 1'b1;
pika_color[5547] <= 1'b1;
pika_color[5597] <= 1'b1;
pika_color[5598] <= 1'b1;
pika_color[5599] <= 1'b1;
pika_color[5600] <= 1'b1;
pika_color[5601] <= 1'b1;
pika_color[5660] <= 1'b1;
pika_color[5661] <= 1'b1;
pika_color[5662] <= 1'b1;
pika_color[5711] <= 1'b1;
pika_color[5712] <= 1'b1;
pika_color[5716] <= 1'b1;
pika_color[5776] <= 1'b1;
pika_color[5777] <= 1'b1;
pika_color[5826] <= 1'b1;
pika_color[5831] <= 1'b1;
pika_color[5832] <= 1'b1;
pika_color[5892] <= 1'b1;
pika_color[5941] <= 1'b1;
pika_color[5947] <= 1'b1;
pika_color[5948] <= 1'b1;
pika_color[6007] <= 1'b1;
pika_color[6044] <= 1'b1;
pika_color[6045] <= 1'b1;
pika_color[6046] <= 1'b1;
pika_color[6047] <= 1'b1;
pika_color[6056] <= 1'b1;
pika_color[6063] <= 1'b1;
pika_color[6122] <= 1'b1;
pika_color[6157] <= 1'b1;
pika_color[6158] <= 1'b1;
pika_color[6159] <= 1'b1;
pika_color[6170] <= 1'b1;
pika_color[6171] <= 1'b1;
pika_color[6178] <= 1'b1;
pika_color[6179] <= 1'b1;
pika_color[6237] <= 1'b1;
pika_color[6285] <= 1'b1;
pika_color[6294] <= 1'b1;
pika_color[6353] <= 1'b1;
pika_color[6400] <= 1'b1;
pika_color[6409] <= 1'b1;
pika_color[6410] <= 1'b1;
pika_color[6468] <= 1'b1;
pika_color[6515] <= 1'b1;
pika_color[6525] <= 1'b1;
pika_color[6583] <= 1'b1;
pika_color[6630] <= 1'b1;
pika_color[6640] <= 1'b1;
pika_color[6698] <= 1'b1;
pika_color[6709] <= 1'b1;
pika_color[6710] <= 1'b1;
pika_color[6711] <= 1'b1;
pika_color[6712] <= 1'b1;
pika_color[6713] <= 1'b1;
pika_color[6714] <= 1'b1;
pika_color[6715] <= 1'b1;
pika_color[6745] <= 1'b1;
pika_color[6755] <= 1'b1;
pika_color[6813] <= 1'b1;
pika_color[6839] <= 1'b1;
pika_color[6840] <= 1'b1;
pika_color[6841] <= 1'b1;
pika_color[6860] <= 1'b1;
pika_color[6870] <= 1'b1;
pika_color[6871] <= 1'b1;
pika_color[6928] <= 1'b1;
pika_color[6952] <= 1'b1;
pika_color[6953] <= 1'b1;
pika_color[6954] <= 1'b1;
pika_color[6955] <= 1'b1;
pika_color[6956] <= 1'b1;
pika_color[6975] <= 1'b1;
pika_color[6986] <= 1'b1;
pika_color[7043] <= 1'b1;
pika_color[7044] <= 1'b1;
pika_color[7068] <= 1'b1;
pika_color[7069] <= 1'b1;
pika_color[7070] <= 1'b1;
pika_color[7090] <= 1'b1;
pika_color[7101] <= 1'b1;
pika_color[7159] <= 1'b1;
pika_color[7205] <= 1'b1;
pika_color[7216] <= 1'b1;
pika_color[7274] <= 1'b1;
pika_color[7320] <= 1'b1;
pika_color[7331] <= 1'b1;
pika_color[7389] <= 1'b1;
pika_color[7435] <= 1'b1;
pika_color[7446] <= 1'b1;
pika_color[7504] <= 1'b1;
pika_color[7530] <= 1'b1;
pika_color[7531] <= 1'b1;
pika_color[7532] <= 1'b1;
pika_color[7533] <= 1'b1;
pika_color[7534] <= 1'b1;
pika_color[7535] <= 1'b1;
pika_color[7536] <= 1'b1;
pika_color[7550] <= 1'b1;
pika_color[7561] <= 1'b1;
pika_color[7619] <= 1'b1;
pika_color[7643] <= 1'b1;
pika_color[7644] <= 1'b1;
pika_color[7645] <= 1'b1;
pika_color[7651] <= 1'b1;
pika_color[7665] <= 1'b1;
pika_color[7676] <= 1'b1;
pika_color[7734] <= 1'b1;
pika_color[7756] <= 1'b1;
pika_color[7757] <= 1'b1;
pika_color[7758] <= 1'b1;
pika_color[7766] <= 1'b1;
pika_color[7780] <= 1'b1;
pika_color[7791] <= 1'b1;
pika_color[7792] <= 1'b1;
pika_color[7849] <= 1'b1;
pika_color[7850] <= 1'b1;
pika_color[7870] <= 1'b1;
pika_color[7871] <= 1'b1;
pika_color[7876] <= 1'b1;
pika_color[7877] <= 1'b1;
pika_color[7878] <= 1'b1;
pika_color[7879] <= 1'b1;
pika_color[7880] <= 1'b1;
pika_color[7881] <= 1'b1;
pika_color[7895] <= 1'b1;
pika_color[7907] <= 1'b1;
pika_color[7965] <= 1'b1;
pika_color[7985] <= 1'b1;
pika_color[7986] <= 1'b1;
pika_color[7989] <= 1'b1;
pika_color[7990] <= 1'b1;
pika_color[7991] <= 1'b1;
pika_color[7996] <= 1'b1;
pika_color[8010] <= 1'b1;
pika_color[8022] <= 1'b1;
pika_color[8080] <= 1'b1;
pika_color[8101] <= 1'b1;
pika_color[8103] <= 1'b1;
pika_color[8104] <= 1'b1;
pika_color[8110] <= 1'b1;
pika_color[8111] <= 1'b1;
pika_color[8125] <= 1'b1;
pika_color[8137] <= 1'b1;
pika_color[8195] <= 1'b1;
pika_color[8196] <= 1'b1;
pika_color[8216] <= 1'b1;
pika_color[8217] <= 1'b1;
pika_color[8218] <= 1'b1;
pika_color[8224] <= 1'b1;
pika_color[8225] <= 1'b1;
pika_color[8240] <= 1'b1;
pika_color[8252] <= 1'b1;
pika_color[8311] <= 1'b1;
pika_color[8312] <= 1'b1;
pika_color[8332] <= 1'b1;
pika_color[8333] <= 1'b1;
pika_color[8334] <= 1'b1;
pika_color[8338] <= 1'b1;
pika_color[8339] <= 1'b1;
pika_color[8354] <= 1'b1;
pika_color[8355] <= 1'b1;
pika_color[8367] <= 1'b1;
pika_color[8426] <= 1'b1;
pika_color[8427] <= 1'b1;
pika_color[8428] <= 1'b1;
pika_color[8449] <= 1'b1;
pika_color[8450] <= 1'b1;
pika_color[8451] <= 1'b1;
pika_color[8452] <= 1'b1;
pika_color[8453] <= 1'b1;
pika_color[8469] <= 1'b1;
pika_color[8482] <= 1'b1;
pika_color[8541] <= 1'b1;
pika_color[8543] <= 1'b1;
pika_color[8544] <= 1'b1;
pika_color[8545] <= 1'b1;
pika_color[8583] <= 1'b1;
pika_color[8584] <= 1'b1;
pika_color[8597] <= 1'b1;
pika_color[8656] <= 1'b1;
pika_color[8660] <= 1'b1;
pika_color[8661] <= 1'b1;
pika_color[8698] <= 1'b1;
pika_color[8712] <= 1'b1;
pika_color[8770] <= 1'b1;
pika_color[8776] <= 1'b1;
pika_color[8777] <= 1'b1;
pika_color[8778] <= 1'b1;
pika_color[8812] <= 1'b1;
pika_color[8827] <= 1'b1;
pika_color[8885] <= 1'b1;
pika_color[8893] <= 1'b1;
pika_color[8894] <= 1'b1;
pika_color[8927] <= 1'b1;
pika_color[8942] <= 1'b1;
pika_color[8999] <= 1'b1;
pika_color[9009] <= 1'b1;
pika_color[9010] <= 1'b1;
pika_color[9057] <= 1'b1;
pika_color[9114] <= 1'b1;
pika_color[9172] <= 1'b1;
pika_color[9228] <= 1'b1;
pika_color[9229] <= 1'b1;
pika_color[9287] <= 1'b1;
pika_color[9343] <= 1'b1;
pika_color[9402] <= 1'b1;
pika_color[9458] <= 1'b1;
pika_color[9517] <= 1'b1;
pika_color[9573] <= 1'b1;
pika_color[9632] <= 1'b1;
pika_color[9687] <= 1'b1;
pika_color[9688] <= 1'b1;
pika_color[9747] <= 1'b1;
pika_color[9802] <= 1'b1;
pika_color[9862] <= 1'b1;
pika_color[9917] <= 1'b1;
pika_color[9977] <= 1'b1;
pika_color[10032] <= 1'b1;
pika_color[10092] <= 1'b1;
pika_color[10147] <= 1'b1;
pika_color[10148] <= 1'b1;
pika_color[10168] <= 1'b1;
pika_color[10169] <= 1'b1;
pika_color[10170] <= 1'b1;
pika_color[10171] <= 1'b1;
pika_color[10172] <= 1'b1;
pika_color[10173] <= 1'b1;
pika_color[10174] <= 1'b1;
pika_color[10207] <= 1'b1;
pika_color[10263] <= 1'b1;
pika_color[10282] <= 1'b1;
pika_color[10283] <= 1'b1;
pika_color[10322] <= 1'b1;
pika_color[10378] <= 1'b1;
pika_color[10397] <= 1'b1;
pika_color[10437] <= 1'b1;
pika_color[10493] <= 1'b1;
pika_color[10494] <= 1'b1;
pika_color[10512] <= 1'b1;
pika_color[10552] <= 1'b1;
pika_color[10609] <= 1'b1;
pika_color[10627] <= 1'b1;
pika_color[10628] <= 1'b1;
pika_color[10667] <= 1'b1;
pika_color[10724] <= 1'b1;
pika_color[10743] <= 1'b1;
pika_color[10782] <= 1'b1;
pika_color[10840] <= 1'b1;
pika_color[10858] <= 1'b1;
pika_color[10859] <= 1'b1;
pika_color[10897] <= 1'b1;
pika_color[10955] <= 1'b1;
pika_color[10956] <= 1'b1;
pika_color[10974] <= 1'b1;
pika_color[11012] <= 1'b1;
pika_color[11070] <= 1'b1;
pika_color[11071] <= 1'b1;
pika_color[11072] <= 1'b1;
pika_color[11089] <= 1'b1;
pika_color[11127] <= 1'b1;
pika_color[11185] <= 1'b1;
pika_color[11187] <= 1'b1;
pika_color[11204] <= 1'b1;
pika_color[11242] <= 1'b1;
pika_color[11300] <= 1'b1;
pika_color[11302] <= 1'b1;
pika_color[11303] <= 1'b1;
pika_color[11319] <= 1'b1;
pika_color[11357] <= 1'b1;
pika_color[11414] <= 1'b1;
pika_color[11415] <= 1'b1;
pika_color[11418] <= 1'b1;
pika_color[11419] <= 1'b1;
pika_color[11434] <= 1'b1;
pika_color[11472] <= 1'b1;
pika_color[11473] <= 1'b1;
pika_color[11529] <= 1'b1;
pika_color[11534] <= 1'b1;
pika_color[11535] <= 1'b1;
pika_color[11548] <= 1'b1;
pika_color[11549] <= 1'b1;
pika_color[11588] <= 1'b1;
pika_color[11644] <= 1'b1;
pika_color[11650] <= 1'b1;
pika_color[11651] <= 1'b1;
pika_color[11663] <= 1'b1;
pika_color[11703] <= 1'b1;
pika_color[11759] <= 1'b1;
pika_color[11766] <= 1'b1;
pika_color[11767] <= 1'b1;
pika_color[11768] <= 1'b1;
pika_color[11778] <= 1'b1;
pika_color[11818] <= 1'b1;
pika_color[11873] <= 1'b1;
pika_color[11883] <= 1'b1;
pika_color[11884] <= 1'b1;
pika_color[11892] <= 1'b1;
pika_color[11933] <= 1'b1;
pika_color[11988] <= 1'b1;
pika_color[11999] <= 1'b1;
pika_color[12000] <= 1'b1;
pika_color[12006] <= 1'b1;
pika_color[12007] <= 1'b1;
pika_color[12048] <= 1'b1;
pika_color[12103] <= 1'b1;
pika_color[12115] <= 1'b1;
pika_color[12116] <= 1'b1;
pika_color[12117] <= 1'b1;
pika_color[12119] <= 1'b1;
pika_color[12120] <= 1'b1;
pika_color[12163] <= 1'b1;
pika_color[12218] <= 1'b1;
pika_color[12232] <= 1'b1;
pika_color[12233] <= 1'b1;
pika_color[12234] <= 1'b1;
pika_color[12278] <= 1'b1;
pika_color[12333] <= 1'b1;
pika_color[12393] <= 1'b1;
pika_color[12448] <= 1'b1;
pika_color[12508] <= 1'b1;
pika_color[12563] <= 1'b1;
pika_color[12623] <= 1'b1;
pika_color[12678] <= 1'b1;
pika_color[12738] <= 1'b1;
pika_color[12793] <= 1'b1;
pika_color[12853] <= 1'b1;
pika_color[12908] <= 1'b1;
pika_color[12968] <= 1'b1;
pika_color[13023] <= 1'b1;
pika_color[13083] <= 1'b1;
pika_color[13138] <= 1'b1;
pika_color[13198] <= 1'b1;
pika_color[13253] <= 1'b1;
pika_color[13254] <= 1'b1;
pika_color[13313] <= 1'b1;
pika_color[13369] <= 1'b1;
pika_color[13427] <= 1'b1;
pika_color[13428] <= 1'b1;
pika_color[13484] <= 1'b1;
pika_color[13542] <= 1'b1;
pika_color[13599] <= 1'b1;
pika_color[13600] <= 1'b1;
pika_color[13657] <= 1'b1;
pika_color[13715] <= 1'b1;
pika_color[13772] <= 1'b1;
pika_color[13830] <= 1'b1;
pika_color[13886] <= 1'b1;
pika_color[13887] <= 1'b1;
pika_color[13945] <= 1'b1;
pika_color[13946] <= 1'b1;
pika_color[14001] <= 1'b1;
pika_color[14061] <= 1'b1;
pika_color[14115] <= 1'b1;
pika_color[14116] <= 1'b1;
pika_color[14176] <= 1'b1;
pika_color[14177] <= 1'b1;
pika_color[14230] <= 1'b1;
pika_color[14292] <= 1'b1;
pika_color[14344] <= 1'b1;
pika_color[14345] <= 1'b1;
pika_color[14407] <= 1'b1;
pika_color[14408] <= 1'b1;
pika_color[14458] <= 1'b1;
pika_color[14459] <= 1'b1;
pika_color[14523] <= 1'b1;
pika_color[14524] <= 1'b1;
pika_color[14547] <= 1'b1;
pika_color[14548] <= 1'b1;
pika_color[14549] <= 1'b1;
pika_color[14550] <= 1'b1;
pika_color[14551] <= 1'b1;
pika_color[14552] <= 1'b1;
pika_color[14572] <= 1'b1;
pika_color[14573] <= 1'b1;
pika_color[14639] <= 1'b1;
pika_color[14640] <= 1'b1;
pika_color[14654] <= 1'b1;
pika_color[14655] <= 1'b1;
pika_color[14656] <= 1'b1;
pika_color[14657] <= 1'b1;
pika_color[14658] <= 1'b1;
pika_color[14659] <= 1'b1;
pika_color[14660] <= 1'b1;
pika_color[14661] <= 1'b1;
pika_color[14662] <= 1'b1;
pika_color[14667] <= 1'b1;
pika_color[14668] <= 1'b1;
pika_color[14669] <= 1'b1;
pika_color[14685] <= 1'b1;
pika_color[14686] <= 1'b1;
pika_color[14687] <= 1'b1;
pika_color[14755] <= 1'b1;
pika_color[14756] <= 1'b1;
pika_color[14757] <= 1'b1;
pika_color[14758] <= 1'b1;
pika_color[14768] <= 1'b1;
pika_color[14784] <= 1'b1;
pika_color[14785] <= 1'b1;
pika_color[14786] <= 1'b1;
pika_color[14787] <= 1'b1;
pika_color[14788] <= 1'b1;
pika_color[14789] <= 1'b1;
pika_color[14799] <= 1'b1;
pika_color[14800] <= 1'b1;
pika_color[14873] <= 1'b1;
pika_color[14874] <= 1'b1;
pika_color[14883] <= 1'b1;
pika_color[14904] <= 1'b1;
pika_color[14905] <= 1'b1;
pika_color[14906] <= 1'b1;
pika_color[14913] <= 1'b1;
pika_color[14914] <= 1'b1;
pika_color[14989] <= 1'b1;
pika_color[14990] <= 1'b1;
pika_color[14991] <= 1'b1;
pika_color[14992] <= 1'b1;
pika_color[14998] <= 1'b1;
pika_color[15021] <= 1'b1;
pika_color[15028] <= 1'b1;
pika_color[15106] <= 1'b1;
pika_color[15107] <= 1'b1;
pika_color[15113] <= 1'b1;
pika_color[15114] <= 1'b1;
pika_color[15136] <= 1'b1;
pika_color[15143] <= 1'b1;
pika_color[15144] <= 1'b1;
pika_color[15221] <= 1'b1;
pika_color[15229] <= 1'b1;
pika_color[15230] <= 1'b1;
pika_color[15250] <= 1'b1;
pika_color[15251] <= 1'b1;
pika_color[15259] <= 1'b1;
pika_color[15260] <= 1'b1;
pika_color[15336] <= 1'b1;
pika_color[15345] <= 1'b1;
pika_color[15365] <= 1'b1;
pika_color[15375] <= 1'b1;
pika_color[15450] <= 1'b1;
pika_color[15451] <= 1'b1;
pika_color[15461] <= 1'b1;
pika_color[15480] <= 1'b1;
pika_color[15490] <= 1'b1;
pika_color[15565] <= 1'b1;
pika_color[15576] <= 1'b1;
pika_color[15595] <= 1'b1;
pika_color[15596] <= 1'b1;
pika_color[15597] <= 1'b1;
pika_color[15603] <= 1'b1;
pika_color[15604] <= 1'b1;
pika_color[15605] <= 1'b1;
pika_color[15680] <= 1'b1;
pika_color[15681] <= 1'b1;
pika_color[15690] <= 1'b1;
pika_color[15691] <= 1'b1;
pika_color[15713] <= 1'b1;
pika_color[15714] <= 1'b1;
pika_color[15715] <= 1'b1;
pika_color[15716] <= 1'b1;
pika_color[15717] <= 1'b1;
pika_color[15718] <= 1'b1;
pika_color[15796] <= 1'b1;
pika_color[15797] <= 1'b1;
pika_color[15802] <= 1'b1;
pika_color[15803] <= 1'b1;
pika_color[15804] <= 1'b1;
pika_color[15805] <= 1'b1;
pika_color[15912] <= 1'b1;
pika_color[15913] <= 1'b1;
pika_color[15914] <= 1'b1;
pika_color[15915] <= 1'b1;
pika_color[15916] <= 1'b1;
pika_color[15917] <= 1'b1;

		end
		move60, move61, move62, move63, move64, move65, move66, move67, move68, move69:
		begin
		pika_color[820] <= 1'b1;
pika_color[821] <= 1'b1;
pika_color[822] <= 1'b1;
pika_color[930] <= 1'b1;
pika_color[931] <= 1'b1;
pika_color[932] <= 1'b1;
pika_color[935] <= 1'b1;
pika_color[937] <= 1'b1;
pika_color[938] <= 1'b1;
pika_color[939] <= 1'b1;
pika_color[1008] <= 1'b1;
pika_color[1009] <= 1'b1;
pika_color[1010] <= 1'b1;
pika_color[1044] <= 1'b1;
pika_color[1045] <= 1'b1;
pika_color[1046] <= 1'b1;
pika_color[1047] <= 1'b1;
pika_color[1048] <= 1'b1;
pika_color[1049] <= 1'b1;
pika_color[1050] <= 1'b1;
pika_color[1054] <= 1'b1;
pika_color[1055] <= 1'b1;
pika_color[1120] <= 1'b1;
pika_color[1121] <= 1'b1;
pika_color[1122] <= 1'b1;
pika_color[1123] <= 1'b1;
pika_color[1124] <= 1'b1;
pika_color[1125] <= 1'b1;
pika_color[1126] <= 1'b1;
pika_color[1127] <= 1'b1;
pika_color[1159] <= 1'b1;
pika_color[1160] <= 1'b1;
pika_color[1161] <= 1'b1;
pika_color[1162] <= 1'b1;
pika_color[1163] <= 1'b1;
pika_color[1164] <= 1'b1;
pika_color[1165] <= 1'b1;
pika_color[1166] <= 1'b1;
pika_color[1167] <= 1'b1;
pika_color[1170] <= 1'b1;
pika_color[1171] <= 1'b1;
pika_color[1231] <= 1'b1;
pika_color[1232] <= 1'b1;
pika_color[1233] <= 1'b1;
pika_color[1234] <= 1'b1;
pika_color[1235] <= 1'b1;
pika_color[1236] <= 1'b1;
pika_color[1237] <= 1'b1;
pika_color[1238] <= 1'b1;
pika_color[1239] <= 1'b1;
pika_color[1240] <= 1'b1;
pika_color[1241] <= 1'b1;
pika_color[1242] <= 1'b1;
pika_color[1243] <= 1'b1;
pika_color[1274] <= 1'b1;
pika_color[1275] <= 1'b1;
pika_color[1276] <= 1'b1;
pika_color[1277] <= 1'b1;
pika_color[1278] <= 1'b1;
pika_color[1279] <= 1'b1;
pika_color[1282] <= 1'b1;
pika_color[1283] <= 1'b1;
pika_color[1284] <= 1'b1;
pika_color[1286] <= 1'b1;
pika_color[1287] <= 1'b1;
pika_color[1344] <= 1'b1;
pika_color[1345] <= 1'b1;
pika_color[1346] <= 1'b1;
pika_color[1351] <= 1'b1;
pika_color[1352] <= 1'b1;
pika_color[1353] <= 1'b1;
pika_color[1354] <= 1'b1;
pika_color[1355] <= 1'b1;
pika_color[1356] <= 1'b1;
pika_color[1357] <= 1'b1;
pika_color[1358] <= 1'b1;
pika_color[1389] <= 1'b1;
pika_color[1390] <= 1'b1;
pika_color[1391] <= 1'b1;
pika_color[1392] <= 1'b1;
pika_color[1393] <= 1'b1;
pika_color[1394] <= 1'b1;
pika_color[1399] <= 1'b1;
pika_color[1400] <= 1'b1;
pika_color[1402] <= 1'b1;
pika_color[1403] <= 1'b1;
pika_color[1457] <= 1'b1;
pika_color[1458] <= 1'b1;
pika_color[1459] <= 1'b1;
pika_color[1466] <= 1'b1;
pika_color[1467] <= 1'b1;
pika_color[1468] <= 1'b1;
pika_color[1469] <= 1'b1;
pika_color[1470] <= 1'b1;
pika_color[1471] <= 1'b1;
pika_color[1472] <= 1'b1;
pika_color[1473] <= 1'b1;
pika_color[1504] <= 1'b1;
pika_color[1505] <= 1'b1;
pika_color[1506] <= 1'b1;
pika_color[1507] <= 1'b1;
pika_color[1508] <= 1'b1;
pika_color[1509] <= 1'b1;
pika_color[1515] <= 1'b1;
pika_color[1516] <= 1'b1;
pika_color[1518] <= 1'b1;
pika_color[1519] <= 1'b1;
pika_color[1570] <= 1'b1;
pika_color[1571] <= 1'b1;
pika_color[1572] <= 1'b1;
pika_color[1580] <= 1'b1;
pika_color[1581] <= 1'b1;
pika_color[1582] <= 1'b1;
pika_color[1583] <= 1'b1;
pika_color[1584] <= 1'b1;
pika_color[1585] <= 1'b1;
pika_color[1586] <= 1'b1;
pika_color[1587] <= 1'b1;
pika_color[1619] <= 1'b1;
pika_color[1620] <= 1'b1;
pika_color[1621] <= 1'b1;
pika_color[1622] <= 1'b1;
pika_color[1623] <= 1'b1;
pika_color[1624] <= 1'b1;
pika_color[1631] <= 1'b1;
pika_color[1632] <= 1'b1;
pika_color[1634] <= 1'b1;
pika_color[1635] <= 1'b1;
pika_color[1684] <= 1'b1;
pika_color[1685] <= 1'b1;
pika_color[1695] <= 1'b1;
pika_color[1696] <= 1'b1;
pika_color[1697] <= 1'b1;
pika_color[1698] <= 1'b1;
pika_color[1699] <= 1'b1;
pika_color[1700] <= 1'b1;
pika_color[1701] <= 1'b1;
pika_color[1702] <= 1'b1;
pika_color[1735] <= 1'b1;
pika_color[1736] <= 1'b1;
pika_color[1737] <= 1'b1;
pika_color[1738] <= 1'b1;
pika_color[1739] <= 1'b1;
pika_color[1747] <= 1'b1;
pika_color[1748] <= 1'b1;
pika_color[1750] <= 1'b1;
pika_color[1798] <= 1'b1;
pika_color[1799] <= 1'b1;
pika_color[1810] <= 1'b1;
pika_color[1811] <= 1'b1;
pika_color[1812] <= 1'b1;
pika_color[1813] <= 1'b1;
pika_color[1814] <= 1'b1;
pika_color[1815] <= 1'b1;
pika_color[1816] <= 1'b1;
pika_color[1850] <= 1'b1;
pika_color[1851] <= 1'b1;
pika_color[1852] <= 1'b1;
pika_color[1853] <= 1'b1;
pika_color[1854] <= 1'b1;
pika_color[1863] <= 1'b1;
pika_color[1864] <= 1'b1;
pika_color[1865] <= 1'b1;
pika_color[1866] <= 1'b1;
pika_color[1912] <= 1'b1;
pika_color[1913] <= 1'b1;
pika_color[1925] <= 1'b1;
pika_color[1926] <= 1'b1;
pika_color[1927] <= 1'b1;
pika_color[1928] <= 1'b1;
pika_color[1929] <= 1'b1;
pika_color[1930] <= 1'b1;
pika_color[1931] <= 1'b1;
pika_color[1966] <= 1'b1;
pika_color[1967] <= 1'b1;
pika_color[1968] <= 1'b1;
pika_color[1979] <= 1'b1;
pika_color[1980] <= 1'b1;
pika_color[1981] <= 1'b1;
pika_color[1982] <= 1'b1;
pika_color[2026] <= 1'b1;
pika_color[2027] <= 1'b1;
pika_color[2039] <= 1'b1;
pika_color[2040] <= 1'b1;
pika_color[2041] <= 1'b1;
pika_color[2042] <= 1'b1;
pika_color[2043] <= 1'b1;
pika_color[2044] <= 1'b1;
pika_color[2045] <= 1'b1;
pika_color[2081] <= 1'b1;
pika_color[2082] <= 1'b1;
pika_color[2083] <= 1'b1;
pika_color[2095] <= 1'b1;
pika_color[2097] <= 1'b1;
pika_color[2098] <= 1'b1;
pika_color[2140] <= 1'b1;
pika_color[2141] <= 1'b1;
pika_color[2154] <= 1'b1;
pika_color[2155] <= 1'b1;
pika_color[2156] <= 1'b1;
pika_color[2157] <= 1'b1;
pika_color[2158] <= 1'b1;
pika_color[2159] <= 1'b1;
pika_color[2197] <= 1'b1;
pika_color[2198] <= 1'b1;
pika_color[2211] <= 1'b1;
pika_color[2213] <= 1'b1;
pika_color[2214] <= 1'b1;
pika_color[2254] <= 1'b1;
pika_color[2255] <= 1'b1;
pika_color[2269] <= 1'b1;
pika_color[2270] <= 1'b1;
pika_color[2271] <= 1'b1;
pika_color[2272] <= 1'b1;
pika_color[2273] <= 1'b1;
pika_color[2274] <= 1'b1;
pika_color[2313] <= 1'b1;
pika_color[2326] <= 1'b1;
pika_color[2327] <= 1'b1;
pika_color[2328] <= 1'b1;
pika_color[2329] <= 1'b1;
pika_color[2330] <= 1'b1;
pika_color[2369] <= 1'b1;
pika_color[2384] <= 1'b1;
pika_color[2385] <= 1'b1;
pika_color[2386] <= 1'b1;
pika_color[2387] <= 1'b1;
pika_color[2388] <= 1'b1;
pika_color[2428] <= 1'b1;
pika_color[2429] <= 1'b1;
pika_color[2442] <= 1'b1;
pika_color[2443] <= 1'b1;
pika_color[2444] <= 1'b1;
pika_color[2445] <= 1'b1;
pika_color[2446] <= 1'b1;
pika_color[2483] <= 1'b1;
pika_color[2484] <= 1'b1;
pika_color[2500] <= 1'b1;
pika_color[2501] <= 1'b1;
pika_color[2502] <= 1'b1;
pika_color[2544] <= 1'b1;
pika_color[2558] <= 1'b1;
pika_color[2559] <= 1'b1;
pika_color[2560] <= 1'b1;
pika_color[2561] <= 1'b1;
pika_color[2597] <= 1'b1;
pika_color[2598] <= 1'b1;
pika_color[2615] <= 1'b1;
pika_color[2616] <= 1'b1;
pika_color[2617] <= 1'b1;
pika_color[2659] <= 1'b1;
pika_color[2660] <= 1'b1;
pika_color[2674] <= 1'b1;
pika_color[2675] <= 1'b1;
pika_color[2676] <= 1'b1;
pika_color[2677] <= 1'b1;
pika_color[2711] <= 1'b1;
pika_color[2712] <= 1'b1;
pika_color[2730] <= 1'b1;
pika_color[2731] <= 1'b1;
pika_color[2775] <= 1'b1;
pika_color[2790] <= 1'b1;
pika_color[2791] <= 1'b1;
pika_color[2792] <= 1'b1;
pika_color[2793] <= 1'b1;
pika_color[2825] <= 1'b1;
pika_color[2826] <= 1'b1;
pika_color[2844] <= 1'b1;
pika_color[2845] <= 1'b1;
pika_color[2890] <= 1'b1;
pika_color[2891] <= 1'b1;
pika_color[2905] <= 1'b1;
pika_color[2906] <= 1'b1;
pika_color[2907] <= 1'b1;
pika_color[2908] <= 1'b1;
pika_color[2917] <= 1'b1;
pika_color[2918] <= 1'b1;
pika_color[2919] <= 1'b1;
pika_color[2920] <= 1'b1;
pika_color[2921] <= 1'b1;
pika_color[2922] <= 1'b1;
pika_color[2923] <= 1'b1;
pika_color[2924] <= 1'b1;
pika_color[2925] <= 1'b1;
pika_color[2926] <= 1'b1;
pika_color[2927] <= 1'b1;
pika_color[2928] <= 1'b1;
pika_color[2939] <= 1'b1;
pika_color[2940] <= 1'b1;
pika_color[2958] <= 1'b1;
pika_color[2959] <= 1'b1;
pika_color[3006] <= 1'b1;
pika_color[3021] <= 1'b1;
pika_color[3022] <= 1'b1;
pika_color[3023] <= 1'b1;
pika_color[3024] <= 1'b1;
pika_color[3028] <= 1'b1;
pika_color[3029] <= 1'b1;
pika_color[3030] <= 1'b1;
pika_color[3031] <= 1'b1;
pika_color[3032] <= 1'b1;
pika_color[3043] <= 1'b1;
pika_color[3044] <= 1'b1;
pika_color[3045] <= 1'b1;
pika_color[3046] <= 1'b1;
pika_color[3047] <= 1'b1;
pika_color[3054] <= 1'b1;
pika_color[3072] <= 1'b1;
pika_color[3073] <= 1'b1;
pika_color[3122] <= 1'b1;
pika_color[3137] <= 1'b1;
pika_color[3138] <= 1'b1;
pika_color[3139] <= 1'b1;
pika_color[3140] <= 1'b1;
pika_color[3141] <= 1'b1;
pika_color[3142] <= 1'b1;
pika_color[3143] <= 1'b1;
pika_color[3162] <= 1'b1;
pika_color[3163] <= 1'b1;
pika_color[3164] <= 1'b1;
pika_color[3165] <= 1'b1;
pika_color[3166] <= 1'b1;
pika_color[3167] <= 1'b1;
pika_color[3168] <= 1'b1;
pika_color[3185] <= 1'b1;
pika_color[3186] <= 1'b1;
pika_color[3187] <= 1'b1;
pika_color[3237] <= 1'b1;
pika_color[3238] <= 1'b1;
pika_color[3253] <= 1'b1;
pika_color[3281] <= 1'b1;
pika_color[3282] <= 1'b1;
pika_color[3299] <= 1'b1;
pika_color[3300] <= 1'b1;
pika_color[3352] <= 1'b1;
pika_color[3353] <= 1'b1;
pika_color[3354] <= 1'b1;
pika_color[3368] <= 1'b1;
pika_color[3369] <= 1'b1;
pika_color[3413] <= 1'b1;
pika_color[3414] <= 1'b1;
pika_color[3467] <= 1'b1;
pika_color[3469] <= 1'b1;
pika_color[3470] <= 1'b1;
pika_color[3484] <= 1'b1;
pika_color[3526] <= 1'b1;
pika_color[3527] <= 1'b1;
pika_color[3528] <= 1'b1;
pika_color[3582] <= 1'b1;
pika_color[3585] <= 1'b1;
pika_color[3640] <= 1'b1;
pika_color[3641] <= 1'b1;
pika_color[3697] <= 1'b1;
pika_color[3700] <= 1'b1;
pika_color[3701] <= 1'b1;
pika_color[3753] <= 1'b1;
pika_color[3754] <= 1'b1;
pika_color[3755] <= 1'b1;
pika_color[3812] <= 1'b1;
pika_color[3813] <= 1'b1;
pika_color[3816] <= 1'b1;
pika_color[3817] <= 1'b1;
pika_color[3866] <= 1'b1;
pika_color[3867] <= 1'b1;
pika_color[3868] <= 1'b1;
pika_color[3928] <= 1'b1;
pika_color[3932] <= 1'b1;
pika_color[3933] <= 1'b1;
pika_color[3979] <= 1'b1;
pika_color[3980] <= 1'b1;
pika_color[3981] <= 1'b1;
pika_color[4043] <= 1'b1;
pika_color[4044] <= 1'b1;
pika_color[4048] <= 1'b1;
pika_color[4094] <= 1'b1;
pika_color[4095] <= 1'b1;
pika_color[4158] <= 1'b1;
pika_color[4159] <= 1'b1;
pika_color[4164] <= 1'b1;
pika_color[4210] <= 1'b1;
pika_color[4211] <= 1'b1;
pika_color[4274] <= 1'b1;
pika_color[4279] <= 1'b1;
pika_color[4280] <= 1'b1;
pika_color[4326] <= 1'b1;
pika_color[4327] <= 1'b1;
pika_color[4389] <= 1'b1;
pika_color[4395] <= 1'b1;
pika_color[4396] <= 1'b1;
pika_color[4442] <= 1'b1;
pika_color[4443] <= 1'b1;
pika_color[4504] <= 1'b1;
pika_color[4505] <= 1'b1;
pika_color[4510] <= 1'b1;
pika_color[4511] <= 1'b1;
pika_color[4558] <= 1'b1;
pika_color[4620] <= 1'b1;
pika_color[4625] <= 1'b1;
pika_color[4673] <= 1'b1;
pika_color[4735] <= 1'b1;
pika_color[4736] <= 1'b1;
pika_color[4740] <= 1'b1;
pika_color[4788] <= 1'b1;
pika_color[4851] <= 1'b1;
pika_color[4852] <= 1'b1;
pika_color[4854] <= 1'b1;
pika_color[4855] <= 1'b1;
pika_color[4903] <= 1'b1;
pika_color[4904] <= 1'b1;
pika_color[4967] <= 1'b1;
pika_color[4968] <= 1'b1;
pika_color[4969] <= 1'b1;
pika_color[5019] <= 1'b1;
pika_color[5083] <= 1'b1;
pika_color[5084] <= 1'b1;
pika_color[5134] <= 1'b1;
pika_color[5199] <= 1'b1;
pika_color[5235] <= 1'b1;
pika_color[5236] <= 1'b1;
pika_color[5237] <= 1'b1;
pika_color[5238] <= 1'b1;
pika_color[5249] <= 1'b1;
pika_color[5314] <= 1'b1;
pika_color[5348] <= 1'b1;
pika_color[5349] <= 1'b1;
pika_color[5364] <= 1'b1;
pika_color[5429] <= 1'b1;
pika_color[5479] <= 1'b1;
pika_color[5543] <= 1'b1;
pika_color[5544] <= 1'b1;
pika_color[5553] <= 1'b1;
pika_color[5554] <= 1'b1;
pika_color[5555] <= 1'b1;
pika_color[5556] <= 1'b1;
pika_color[5557] <= 1'b1;
pika_color[5558] <= 1'b1;
pika_color[5559] <= 1'b1;
pika_color[5594] <= 1'b1;
pika_color[5658] <= 1'b1;
pika_color[5709] <= 1'b1;
pika_color[5773] <= 1'b1;
pika_color[5797] <= 1'b1;
pika_color[5798] <= 1'b1;
pika_color[5799] <= 1'b1;
pika_color[5800] <= 1'b1;
pika_color[5824] <= 1'b1;
pika_color[5825] <= 1'b1;
pika_color[5826] <= 1'b1;
pika_color[5888] <= 1'b1;
pika_color[5911] <= 1'b1;
pika_color[5912] <= 1'b1;
pika_color[5913] <= 1'b1;
pika_color[5914] <= 1'b1;
pika_color[5915] <= 1'b1;
pika_color[5937] <= 1'b1;
pika_color[5938] <= 1'b1;
pika_color[5939] <= 1'b1;
pika_color[5942] <= 1'b1;
pika_color[5943] <= 1'b1;
pika_color[5944] <= 1'b1;
pika_color[5945] <= 1'b1;
pika_color[6003] <= 1'b1;
pika_color[6027] <= 1'b1;
pika_color[6028] <= 1'b1;
pika_color[6052] <= 1'b1;
pika_color[6061] <= 1'b1;
pika_color[6118] <= 1'b1;
pika_color[6166] <= 1'b1;
pika_color[6167] <= 1'b1;
pika_color[6177] <= 1'b1;
pika_color[6233] <= 1'b1;
pika_color[6281] <= 1'b1;
pika_color[6292] <= 1'b1;
pika_color[6293] <= 1'b1;
pika_color[6348] <= 1'b1;
pika_color[6396] <= 1'b1;
pika_color[6408] <= 1'b1;
pika_color[6463] <= 1'b1;
pika_color[6486] <= 1'b1;
pika_color[6487] <= 1'b1;
pika_color[6488] <= 1'b1;
pika_color[6489] <= 1'b1;
pika_color[6490] <= 1'b1;
pika_color[6491] <= 1'b1;
pika_color[6492] <= 1'b1;
pika_color[6493] <= 1'b1;
pika_color[6511] <= 1'b1;
pika_color[6523] <= 1'b1;
pika_color[6578] <= 1'b1;
pika_color[6597] <= 1'b1;
pika_color[6598] <= 1'b1;
pika_color[6599] <= 1'b1;
pika_color[6600] <= 1'b1;
pika_color[6601] <= 1'b1;
pika_color[6626] <= 1'b1;
pika_color[6638] <= 1'b1;
pika_color[6693] <= 1'b1;
pika_color[6741] <= 1'b1;
pika_color[6753] <= 1'b1;
pika_color[6808] <= 1'b1;
pika_color[6856] <= 1'b1;
pika_color[6868] <= 1'b1;
pika_color[6923] <= 1'b1;
pika_color[6971] <= 1'b1;
pika_color[6983] <= 1'b1;
pika_color[7038] <= 1'b1;
pika_color[7085] <= 1'b1;
pika_color[7086] <= 1'b1;
pika_color[7098] <= 1'b1;
pika_color[7154] <= 1'b1;
pika_color[7199] <= 1'b1;
pika_color[7200] <= 1'b1;
pika_color[7213] <= 1'b1;
pika_color[7269] <= 1'b1;
pika_color[7270] <= 1'b1;
pika_color[7314] <= 1'b1;
pika_color[7328] <= 1'b1;
pika_color[7385] <= 1'b1;
pika_color[7428] <= 1'b1;
pika_color[7429] <= 1'b1;
pika_color[7443] <= 1'b1;
pika_color[7500] <= 1'b1;
pika_color[7543] <= 1'b1;
pika_color[7558] <= 1'b1;
pika_color[7615] <= 1'b1;
pika_color[7616] <= 1'b1;
pika_color[7657] <= 1'b1;
pika_color[7658] <= 1'b1;
pika_color[7672] <= 1'b1;
pika_color[7673] <= 1'b1;
pika_color[7731] <= 1'b1;
pika_color[7772] <= 1'b1;
pika_color[7787] <= 1'b1;
pika_color[7846] <= 1'b1;
pika_color[7847] <= 1'b1;
pika_color[7886] <= 1'b1;
pika_color[7902] <= 1'b1;
pika_color[7961] <= 1'b1;
pika_color[7962] <= 1'b1;
pika_color[7963] <= 1'b1;
pika_color[8000] <= 1'b1;
pika_color[8001] <= 1'b1;
pika_color[8017] <= 1'b1;
pika_color[8076] <= 1'b1;
pika_color[8078] <= 1'b1;
pika_color[8079] <= 1'b1;
pika_color[8080] <= 1'b1;
pika_color[8114] <= 1'b1;
pika_color[8115] <= 1'b1;
pika_color[8132] <= 1'b1;
pika_color[8190] <= 1'b1;
pika_color[8195] <= 1'b1;
pika_color[8196] <= 1'b1;
pika_color[8197] <= 1'b1;
pika_color[8229] <= 1'b1;
pika_color[8246] <= 1'b1;
pika_color[8247] <= 1'b1;
pika_color[8305] <= 1'b1;
pika_color[8313] <= 1'b1;
pika_color[8314] <= 1'b1;
pika_color[8315] <= 1'b1;
pika_color[8343] <= 1'b1;
pika_color[8344] <= 1'b1;
pika_color[8361] <= 1'b1;
pika_color[8420] <= 1'b1;
pika_color[8457] <= 1'b1;
pika_color[8458] <= 1'b1;
pika_color[8476] <= 1'b1;
pika_color[8535] <= 1'b1;
pika_color[8572] <= 1'b1;
pika_color[8591] <= 1'b1;
pika_color[8649] <= 1'b1;
pika_color[8650] <= 1'b1;
pika_color[8705] <= 1'b1;
pika_color[8706] <= 1'b1;
pika_color[8764] <= 1'b1;
pika_color[8820] <= 1'b1;
pika_color[8879] <= 1'b1;
pika_color[8934] <= 1'b1;
pika_color[8935] <= 1'b1;
pika_color[8994] <= 1'b1;
pika_color[9049] <= 1'b1;
pika_color[9109] <= 1'b1;
pika_color[9164] <= 1'b1;
pika_color[9223] <= 1'b1;
pika_color[9224] <= 1'b1;
pika_color[9279] <= 1'b1;
pika_color[9338] <= 1'b1;
pika_color[9394] <= 1'b1;
pika_color[9453] <= 1'b1;
pika_color[9509] <= 1'b1;
pika_color[9568] <= 1'b1;
pika_color[9624] <= 1'b1;
pika_color[9683] <= 1'b1;
pika_color[9739] <= 1'b1;
pika_color[9798] <= 1'b1;
pika_color[9823] <= 1'b1;
pika_color[9824] <= 1'b1;
pika_color[9825] <= 1'b1;
pika_color[9854] <= 1'b1;
pika_color[9913] <= 1'b1;
pika_color[9936] <= 1'b1;
pika_color[9937] <= 1'b1;
pika_color[9938] <= 1'b1;
pika_color[9969] <= 1'b1;
pika_color[10028] <= 1'b1;
pika_color[10049] <= 1'b1;
pika_color[10050] <= 1'b1;
pika_color[10084] <= 1'b1;
pika_color[10143] <= 1'b1;
pika_color[10163] <= 1'b1;
pika_color[10164] <= 1'b1;
pika_color[10199] <= 1'b1;
pika_color[10258] <= 1'b1;
pika_color[10277] <= 1'b1;
pika_color[10278] <= 1'b1;
pika_color[10314] <= 1'b1;
pika_color[10373] <= 1'b1;
pika_color[10392] <= 1'b1;
pika_color[10429] <= 1'b1;
pika_color[10488] <= 1'b1;
pika_color[10489] <= 1'b1;
pika_color[10507] <= 1'b1;
pika_color[10544] <= 1'b1;
pika_color[10604] <= 1'b1;
pika_color[10622] <= 1'b1;
pika_color[10659] <= 1'b1;
pika_color[10719] <= 1'b1;
pika_color[10737] <= 1'b1;
pika_color[10774] <= 1'b1;
pika_color[10834] <= 1'b1;
pika_color[10835] <= 1'b1;
pika_color[10852] <= 1'b1;
pika_color[10889] <= 1'b1;
pika_color[10949] <= 1'b1;
pika_color[10950] <= 1'b1;
pika_color[10967] <= 1'b1;
pika_color[11004] <= 1'b1;
pika_color[11064] <= 1'b1;
pika_color[11065] <= 1'b1;
pika_color[11082] <= 1'b1;
pika_color[11119] <= 1'b1;
pika_color[11179] <= 1'b1;
pika_color[11181] <= 1'b1;
pika_color[11197] <= 1'b1;
pika_color[11234] <= 1'b1;
pika_color[11294] <= 1'b1;
pika_color[11296] <= 1'b1;
pika_color[11312] <= 1'b1;
pika_color[11349] <= 1'b1;
pika_color[11409] <= 1'b1;
pika_color[11411] <= 1'b1;
pika_color[11412] <= 1'b1;
pika_color[11427] <= 1'b1;
pika_color[11464] <= 1'b1;
pika_color[11465] <= 1'b1;
pika_color[11524] <= 1'b1;
pika_color[11527] <= 1'b1;
pika_color[11528] <= 1'b1;
pika_color[11542] <= 1'b1;
pika_color[11580] <= 1'b1;
pika_color[11639] <= 1'b1;
pika_color[11643] <= 1'b1;
pika_color[11644] <= 1'b1;
pika_color[11656] <= 1'b1;
pika_color[11657] <= 1'b1;
pika_color[11695] <= 1'b1;
pika_color[11754] <= 1'b1;
pika_color[11759] <= 1'b1;
pika_color[11760] <= 1'b1;
pika_color[11769] <= 1'b1;
pika_color[11770] <= 1'b1;
pika_color[11771] <= 1'b1;
pika_color[11810] <= 1'b1;
pika_color[11869] <= 1'b1;
pika_color[11875] <= 1'b1;
pika_color[11876] <= 1'b1;
pika_color[11882] <= 1'b1;
pika_color[11883] <= 1'b1;
pika_color[11884] <= 1'b1;
pika_color[11925] <= 1'b1;
pika_color[11984] <= 1'b1;
pika_color[11991] <= 1'b1;
pika_color[11992] <= 1'b1;
pika_color[11993] <= 1'b1;
pika_color[11994] <= 1'b1;
pika_color[11995] <= 1'b1;
pika_color[11996] <= 1'b1;
pika_color[11997] <= 1'b1;
pika_color[12040] <= 1'b1;
pika_color[12099] <= 1'b1;
pika_color[12155] <= 1'b1;
pika_color[12214] <= 1'b1;
pika_color[12270] <= 1'b1;
pika_color[12329] <= 1'b1;
pika_color[12385] <= 1'b1;
pika_color[12444] <= 1'b1;
pika_color[12499] <= 1'b1;
pika_color[12500] <= 1'b1;
pika_color[12559] <= 1'b1;
pika_color[12614] <= 1'b1;
pika_color[12674] <= 1'b1;
pika_color[12729] <= 1'b1;
pika_color[12789] <= 1'b1;
pika_color[12844] <= 1'b1;
pika_color[12904] <= 1'b1;
pika_color[12905] <= 1'b1;
pika_color[12959] <= 1'b1;
pika_color[13020] <= 1'b1;
pika_color[13074] <= 1'b1;
pika_color[13135] <= 1'b1;
pika_color[13188] <= 1'b1;
pika_color[13189] <= 1'b1;
pika_color[13250] <= 1'b1;
pika_color[13251] <= 1'b1;
pika_color[13303] <= 1'b1;
pika_color[13366] <= 1'b1;
pika_color[13418] <= 1'b1;
pika_color[13481] <= 1'b1;
pika_color[13532] <= 1'b1;
pika_color[13533] <= 1'b1;
pika_color[13596] <= 1'b1;
pika_color[13647] <= 1'b1;
pika_color[13711] <= 1'b1;
pika_color[13712] <= 1'b1;
pika_color[13762] <= 1'b1;
pika_color[13827] <= 1'b1;
pika_color[13877] <= 1'b1;
pika_color[13942] <= 1'b1;
pika_color[13992] <= 1'b1;
pika_color[14057] <= 1'b1;
pika_color[14058] <= 1'b1;
pika_color[14106] <= 1'b1;
pika_color[14107] <= 1'b1;
pika_color[14173] <= 1'b1;
pika_color[14221] <= 1'b1;
pika_color[14288] <= 1'b1;
pika_color[14289] <= 1'b1;
pika_color[14335] <= 1'b1;
pika_color[14336] <= 1'b1;
pika_color[14404] <= 1'b1;
pika_color[14424] <= 1'b1;
pika_color[14425] <= 1'b1;
pika_color[14426] <= 1'b1;
pika_color[14427] <= 1'b1;
pika_color[14428] <= 1'b1;
pika_color[14429] <= 1'b1;
pika_color[14430] <= 1'b1;
pika_color[14431] <= 1'b1;
pika_color[14449] <= 1'b1;
pika_color[14450] <= 1'b1;
pika_color[14519] <= 1'b1;
pika_color[14520] <= 1'b1;
pika_color[14537] <= 1'b1;
pika_color[14538] <= 1'b1;
pika_color[14539] <= 1'b1;
pika_color[14547] <= 1'b1;
pika_color[14548] <= 1'b1;
pika_color[14564] <= 1'b1;
pika_color[14635] <= 1'b1;
pika_color[14636] <= 1'b1;
pika_color[14650] <= 1'b1;
pika_color[14651] <= 1'b1;
pika_color[14663] <= 1'b1;
pika_color[14664] <= 1'b1;
pika_color[14665] <= 1'b1;
pika_color[14678] <= 1'b1;
pika_color[14679] <= 1'b1;
pika_color[14751] <= 1'b1;
pika_color[14752] <= 1'b1;
pika_color[14753] <= 1'b1;
pika_color[14764] <= 1'b1;
pika_color[14765] <= 1'b1;
pika_color[14780] <= 1'b1;
pika_color[14781] <= 1'b1;
pika_color[14792] <= 1'b1;
pika_color[14793] <= 1'b1;
pika_color[14868] <= 1'b1;
pika_color[14869] <= 1'b1;
pika_color[14879] <= 1'b1;
pika_color[14896] <= 1'b1;
pika_color[14906] <= 1'b1;
pika_color[14907] <= 1'b1;
pika_color[14984] <= 1'b1;
pika_color[14985] <= 1'b1;
pika_color[14986] <= 1'b1;
pika_color[14994] <= 1'b1;
pika_color[15011] <= 1'b1;
pika_color[15021] <= 1'b1;
pika_color[15101] <= 1'b1;
pika_color[15102] <= 1'b1;
pika_color[15103] <= 1'b1;
pika_color[15104] <= 1'b1;
pika_color[15109] <= 1'b1;
pika_color[15126] <= 1'b1;
pika_color[15136] <= 1'b1;
pika_color[15219] <= 1'b1;
pika_color[15224] <= 1'b1;
pika_color[15241] <= 1'b1;
pika_color[15251] <= 1'b1;
pika_color[15333] <= 1'b1;
pika_color[15334] <= 1'b1;
pika_color[15339] <= 1'b1;
pika_color[15340] <= 1'b1;
pika_color[15341] <= 1'b1;
pika_color[15357] <= 1'b1;
pika_color[15365] <= 1'b1;
pika_color[15366] <= 1'b1;
pika_color[15448] <= 1'b1;
pika_color[15456] <= 1'b1;
pika_color[15473] <= 1'b1;
pika_color[15474] <= 1'b1;
pika_color[15475] <= 1'b1;
pika_color[15476] <= 1'b1;
pika_color[15477] <= 1'b1;
pika_color[15478] <= 1'b1;
pika_color[15479] <= 1'b1;
pika_color[15480] <= 1'b1;
pika_color[15563] <= 1'b1;
pika_color[15571] <= 1'b1;
pika_color[15678] <= 1'b1;
pika_color[15685] <= 1'b1;
pika_color[15686] <= 1'b1;
pika_color[15793] <= 1'b1;
pika_color[15794] <= 1'b1;
pika_color[15795] <= 1'b1;
pika_color[15796] <= 1'b1;
pika_color[15797] <= 1'b1;
pika_color[15798] <= 1'b1;
pika_color[15799] <= 1'b1;
pika_color[15800] <= 1'b1;

		end
		move70, move71, move72, move73, move74, move75, move76, move77, move78, move79:
begin
pika_color[819] <= 1'b1;
pika_color[820] <= 1'b1;
pika_color[821] <= 1'b1;
pika_color[822] <= 1'b1;
pika_color[823] <= 1'b1;
pika_color[929] <= 1'b1;
pika_color[930] <= 1'b1;
pika_color[931] <= 1'b1;
pika_color[932] <= 1'b1;
pika_color[934] <= 1'b1;
pika_color[935] <= 1'b1;
pika_color[936] <= 1'b1;
pika_color[937] <= 1'b1;
pika_color[938] <= 1'b1;
pika_color[939] <= 1'b1;
pika_color[940] <= 1'b1;
pika_color[941] <= 1'b1;
pika_color[1043] <= 1'b1;
pika_color[1044] <= 1'b1;
pika_color[1047] <= 1'b1;
pika_color[1048] <= 1'b1;
pika_color[1049] <= 1'b1;
pika_color[1050] <= 1'b1;
pika_color[1051] <= 1'b1;
pika_color[1052] <= 1'b1;
pika_color[1053] <= 1'b1;
pika_color[1054] <= 1'b1;
pika_color[1055] <= 1'b1;
pika_color[1056] <= 1'b1;
pika_color[1057] <= 1'b1;
pika_color[1058] <= 1'b1;
pika_color[1158] <= 1'b1;
pika_color[1163] <= 1'b1;
pika_color[1164] <= 1'b1;
pika_color[1165] <= 1'b1;
pika_color[1166] <= 1'b1;
pika_color[1167] <= 1'b1;
pika_color[1168] <= 1'b1;
pika_color[1169] <= 1'b1;
pika_color[1170] <= 1'b1;
pika_color[1173] <= 1'b1;
pika_color[1174] <= 1'b1;
pika_color[1273] <= 1'b1;
pika_color[1279] <= 1'b1;
pika_color[1280] <= 1'b1;
pika_color[1281] <= 1'b1;
pika_color[1282] <= 1'b1;
pika_color[1283] <= 1'b1;
pika_color[1284] <= 1'b1;
pika_color[1289] <= 1'b1;
pika_color[1290] <= 1'b1;
pika_color[1388] <= 1'b1;
pika_color[1394] <= 1'b1;
pika_color[1395] <= 1'b1;
pika_color[1396] <= 1'b1;
pika_color[1397] <= 1'b1;
pika_color[1398] <= 1'b1;
pika_color[1399] <= 1'b1;
pika_color[1405] <= 1'b1;
pika_color[1406] <= 1'b1;
pika_color[1503] <= 1'b1;
pika_color[1509] <= 1'b1;
pika_color[1510] <= 1'b1;
pika_color[1511] <= 1'b1;
pika_color[1512] <= 1'b1;
pika_color[1513] <= 1'b1;
pika_color[1514] <= 1'b1;
pika_color[1521] <= 1'b1;
pika_color[1522] <= 1'b1;
pika_color[1618] <= 1'b1;
pika_color[1624] <= 1'b1;
pika_color[1625] <= 1'b1;
pika_color[1626] <= 1'b1;
pika_color[1627] <= 1'b1;
pika_color[1628] <= 1'b1;
pika_color[1629] <= 1'b1;
pika_color[1637] <= 1'b1;
pika_color[1638] <= 1'b1;
pika_color[1733] <= 1'b1;
pika_color[1740] <= 1'b1;
pika_color[1741] <= 1'b1;
pika_color[1742] <= 1'b1;
pika_color[1743] <= 1'b1;
pika_color[1744] <= 1'b1;
pika_color[1753] <= 1'b1;
pika_color[1754] <= 1'b1;
pika_color[1848] <= 1'b1;
pika_color[1855] <= 1'b1;
pika_color[1856] <= 1'b1;
pika_color[1857] <= 1'b1;
pika_color[1858] <= 1'b1;
pika_color[1859] <= 1'b1;
pika_color[1869] <= 1'b1;
pika_color[1870] <= 1'b1;
pika_color[1963] <= 1'b1;
pika_color[1970] <= 1'b1;
pika_color[1971] <= 1'b1;
pika_color[1972] <= 1'b1;
pika_color[1973] <= 1'b1;
pika_color[1974] <= 1'b1;
pika_color[1985] <= 1'b1;
pika_color[2078] <= 1'b1;
pika_color[2086] <= 1'b1;
pika_color[2087] <= 1'b1;
pika_color[2088] <= 1'b1;
pika_color[2089] <= 1'b1;
pika_color[2100] <= 1'b1;
pika_color[2101] <= 1'b1;
pika_color[2193] <= 1'b1;
pika_color[2201] <= 1'b1;
pika_color[2202] <= 1'b1;
pika_color[2203] <= 1'b1;
pika_color[2204] <= 1'b1;
pika_color[2216] <= 1'b1;
pika_color[2217] <= 1'b1;
pika_color[2308] <= 1'b1;
pika_color[2317] <= 1'b1;
pika_color[2318] <= 1'b1;
pika_color[2319] <= 1'b1;
pika_color[2332] <= 1'b1;
pika_color[2333] <= 1'b1;
pika_color[2423] <= 1'b1;
pika_color[2432] <= 1'b1;
pika_color[2433] <= 1'b1;
pika_color[2448] <= 1'b1;
pika_color[2449] <= 1'b1;
pika_color[2538] <= 1'b1;
pika_color[2539] <= 1'b1;
pika_color[2547] <= 1'b1;
pika_color[2548] <= 1'b1;
pika_color[2564] <= 1'b1;
pika_color[2654] <= 1'b1;
pika_color[2663] <= 1'b1;
pika_color[2679] <= 1'b1;
pika_color[2680] <= 1'b1;
pika_color[2769] <= 1'b1;
pika_color[2778] <= 1'b1;
pika_color[2779] <= 1'b1;
pika_color[2795] <= 1'b1;
pika_color[2884] <= 1'b1;
pika_color[2894] <= 1'b1;
pika_color[2895] <= 1'b1;
pika_color[2911] <= 1'b1;
pika_color[2999] <= 1'b1;
pika_color[3010] <= 1'b1;
pika_color[3026] <= 1'b1;
pika_color[3027] <= 1'b1;
pika_color[3114] <= 1'b1;
pika_color[3126] <= 1'b1;
pika_color[3142] <= 1'b1;
pika_color[3198] <= 1'b1;
pika_color[3199] <= 1'b1;
pika_color[3200] <= 1'b1;
pika_color[3201] <= 1'b1;
pika_color[3202] <= 1'b1;
pika_color[3203] <= 1'b1;
pika_color[3229] <= 1'b1;
pika_color[3241] <= 1'b1;
pika_color[3242] <= 1'b1;
pika_color[3257] <= 1'b1;
pika_color[3258] <= 1'b1;
pika_color[3264] <= 1'b1;
pika_color[3265] <= 1'b1;
pika_color[3266] <= 1'b1;
pika_color[3267] <= 1'b1;
pika_color[3268] <= 1'b1;
pika_color[3269] <= 1'b1;
pika_color[3270] <= 1'b1;
pika_color[3271] <= 1'b1;
pika_color[3272] <= 1'b1;
pika_color[3273] <= 1'b1;
pika_color[3274] <= 1'b1;
pika_color[3275] <= 1'b1;
pika_color[3306] <= 1'b1;
pika_color[3307] <= 1'b1;
pika_color[3308] <= 1'b1;
pika_color[3309] <= 1'b1;
pika_color[3310] <= 1'b1;
pika_color[3311] <= 1'b1;
pika_color[3312] <= 1'b1;
pika_color[3313] <= 1'b1;
pika_color[3319] <= 1'b1;
pika_color[3320] <= 1'b1;
pika_color[3321] <= 1'b1;
pika_color[3322] <= 1'b1;
pika_color[3323] <= 1'b1;
pika_color[3324] <= 1'b1;
pika_color[3344] <= 1'b1;
pika_color[3357] <= 1'b1;
pika_color[3358] <= 1'b1;
pika_color[3373] <= 1'b1;
pika_color[3375] <= 1'b1;
pika_color[3376] <= 1'b1;
pika_color[3377] <= 1'b1;
pika_color[3378] <= 1'b1;
pika_color[3390] <= 1'b1;
pika_color[3391] <= 1'b1;
pika_color[3392] <= 1'b1;
pika_color[3393] <= 1'b1;
pika_color[3394] <= 1'b1;
pika_color[3395] <= 1'b1;
pika_color[3417] <= 1'b1;
pika_color[3418] <= 1'b1;
pika_color[3419] <= 1'b1;
pika_color[3420] <= 1'b1;
pika_color[3421] <= 1'b1;
pika_color[3437] <= 1'b1;
pika_color[3438] <= 1'b1;
pika_color[3439] <= 1'b1;
pika_color[3440] <= 1'b1;
pika_color[3441] <= 1'b1;
pika_color[3459] <= 1'b1;
pika_color[3460] <= 1'b1;
pika_color[3473] <= 1'b1;
pika_color[3488] <= 1'b1;
pika_color[3489] <= 1'b1;
pika_color[3490] <= 1'b1;
pika_color[3510] <= 1'b1;
pika_color[3511] <= 1'b1;
pika_color[3512] <= 1'b1;
pika_color[3513] <= 1'b1;
pika_color[3527] <= 1'b1;
pika_color[3528] <= 1'b1;
pika_color[3529] <= 1'b1;
pika_color[3530] <= 1'b1;
pika_color[3531] <= 1'b1;
pika_color[3532] <= 1'b1;
pika_color[3552] <= 1'b1;
pika_color[3553] <= 1'b1;
pika_color[3554] <= 1'b1;
pika_color[3555] <= 1'b1;
pika_color[3556] <= 1'b1;
pika_color[3557] <= 1'b1;
pika_color[3558] <= 1'b1;
pika_color[3559] <= 1'b1;
pika_color[3575] <= 1'b1;
pika_color[3588] <= 1'b1;
pika_color[3589] <= 1'b1;
pika_color[3603] <= 1'b1;
pika_color[3628] <= 1'b1;
pika_color[3629] <= 1'b1;
pika_color[3639] <= 1'b1;
pika_color[3640] <= 1'b1;
pika_color[3641] <= 1'b1;
pika_color[3642] <= 1'b1;
pika_color[3666] <= 1'b1;
pika_color[3667] <= 1'b1;
pika_color[3668] <= 1'b1;
pika_color[3669] <= 1'b1;
pika_color[3670] <= 1'b1;
pika_color[3671] <= 1'b1;
pika_color[3672] <= 1'b1;
pika_color[3673] <= 1'b1;
pika_color[3674] <= 1'b1;
pika_color[3675] <= 1'b1;
pika_color[3690] <= 1'b1;
pika_color[3704] <= 1'b1;
pika_color[3705] <= 1'b1;
pika_color[3744] <= 1'b1;
pika_color[3745] <= 1'b1;
pika_color[3746] <= 1'b1;
pika_color[3747] <= 1'b1;
pika_color[3750] <= 1'b1;
pika_color[3751] <= 1'b1;
pika_color[3752] <= 1'b1;
pika_color[3753] <= 1'b1;
pika_color[3754] <= 1'b1;
pika_color[3780] <= 1'b1;
pika_color[3781] <= 1'b1;
pika_color[3782] <= 1'b1;
pika_color[3783] <= 1'b1;
pika_color[3784] <= 1'b1;
pika_color[3785] <= 1'b1;
pika_color[3786] <= 1'b1;
pika_color[3787] <= 1'b1;
pika_color[3788] <= 1'b1;
pika_color[3789] <= 1'b1;
pika_color[3790] <= 1'b1;
pika_color[3805] <= 1'b1;
pika_color[3820] <= 1'b1;
pika_color[3821] <= 1'b1;
pika_color[3862] <= 1'b1;
pika_color[3863] <= 1'b1;
pika_color[3864] <= 1'b1;
pika_color[3865] <= 1'b1;
pika_color[3894] <= 1'b1;
pika_color[3895] <= 1'b1;
pika_color[3896] <= 1'b1;
pika_color[3897] <= 1'b1;
pika_color[3898] <= 1'b1;
pika_color[3899] <= 1'b1;
pika_color[3900] <= 1'b1;
pika_color[3901] <= 1'b1;
pika_color[3902] <= 1'b1;
pika_color[3903] <= 1'b1;
pika_color[3904] <= 1'b1;
pika_color[3920] <= 1'b1;
pika_color[3936] <= 1'b1;
pika_color[3937] <= 1'b1;
pika_color[4008] <= 1'b1;
pika_color[4009] <= 1'b1;
pika_color[4010] <= 1'b1;
pika_color[4011] <= 1'b1;
pika_color[4012] <= 1'b1;
pika_color[4013] <= 1'b1;
pika_color[4014] <= 1'b1;
pika_color[4015] <= 1'b1;
pika_color[4016] <= 1'b1;
pika_color[4017] <= 1'b1;
pika_color[4035] <= 1'b1;
pika_color[4052] <= 1'b1;
pika_color[4053] <= 1'b1;
pika_color[4123] <= 1'b1;
pika_color[4124] <= 1'b1;
pika_color[4125] <= 1'b1;
pika_color[4126] <= 1'b1;
pika_color[4127] <= 1'b1;
pika_color[4128] <= 1'b1;
pika_color[4129] <= 1'b1;
pika_color[4130] <= 1'b1;
pika_color[4131] <= 1'b1;
pika_color[4150] <= 1'b1;
pika_color[4151] <= 1'b1;
pika_color[4168] <= 1'b1;
pika_color[4169] <= 1'b1;
pika_color[4237] <= 1'b1;
pika_color[4238] <= 1'b1;
pika_color[4239] <= 1'b1;
pika_color[4240] <= 1'b1;
pika_color[4241] <= 1'b1;
pika_color[4242] <= 1'b1;
pika_color[4243] <= 1'b1;
pika_color[4244] <= 1'b1;
pika_color[4245] <= 1'b1;
pika_color[4266] <= 1'b1;
pika_color[4284] <= 1'b1;
pika_color[4285] <= 1'b1;
pika_color[4351] <= 1'b1;
pika_color[4352] <= 1'b1;
pika_color[4353] <= 1'b1;
pika_color[4354] <= 1'b1;
pika_color[4355] <= 1'b1;
pika_color[4356] <= 1'b1;
pika_color[4357] <= 1'b1;
pika_color[4358] <= 1'b1;
pika_color[4381] <= 1'b1;
pika_color[4400] <= 1'b1;
pika_color[4466] <= 1'b1;
pika_color[4467] <= 1'b1;
pika_color[4468] <= 1'b1;
pika_color[4469] <= 1'b1;
pika_color[4470] <= 1'b1;
pika_color[4471] <= 1'b1;
pika_color[4496] <= 1'b1;
pika_color[4514] <= 1'b1;
pika_color[4515] <= 1'b1;
pika_color[4580] <= 1'b1;
pika_color[4581] <= 1'b1;
pika_color[4582] <= 1'b1;
pika_color[4583] <= 1'b1;
pika_color[4584] <= 1'b1;
pika_color[4611] <= 1'b1;
pika_color[4629] <= 1'b1;
pika_color[4693] <= 1'b1;
pika_color[4694] <= 1'b1;
pika_color[4695] <= 1'b1;
pika_color[4696] <= 1'b1;
pika_color[4726] <= 1'b1;
pika_color[4727] <= 1'b1;
pika_color[4744] <= 1'b1;
pika_color[4787] <= 1'b1;
pika_color[4788] <= 1'b1;
pika_color[4789] <= 1'b1;
pika_color[4797] <= 1'b1;
pika_color[4798] <= 1'b1;
pika_color[4799] <= 1'b1;
pika_color[4800] <= 1'b1;
pika_color[4801] <= 1'b1;
pika_color[4802] <= 1'b1;
pika_color[4803] <= 1'b1;
pika_color[4804] <= 1'b1;
pika_color[4805] <= 1'b1;
pika_color[4806] <= 1'b1;
pika_color[4807] <= 1'b1;
pika_color[4808] <= 1'b1;
pika_color[4842] <= 1'b1;
pika_color[4858] <= 1'b1;
pika_color[4859] <= 1'b1;
pika_color[4904] <= 1'b1;
pika_color[4905] <= 1'b1;
pika_color[4906] <= 1'b1;
pika_color[4907] <= 1'b1;
pika_color[4908] <= 1'b1;
pika_color[4909] <= 1'b1;
pika_color[4910] <= 1'b1;
pika_color[4911] <= 1'b1;
pika_color[4912] <= 1'b1;
pika_color[4957] <= 1'b1;
pika_color[4958] <= 1'b1;
pika_color[4973] <= 1'b1;
pika_color[5020] <= 1'b1;
pika_color[5021] <= 1'b1;
pika_color[5073] <= 1'b1;
pika_color[5074] <= 1'b1;
pika_color[5087] <= 1'b1;
pika_color[5088] <= 1'b1;
pika_color[5136] <= 1'b1;
pika_color[5137] <= 1'b1;
pika_color[5189] <= 1'b1;
pika_color[5190] <= 1'b1;
pika_color[5202] <= 1'b1;
pika_color[5252] <= 1'b1;
pika_color[5305] <= 1'b1;
pika_color[5306] <= 1'b1;
pika_color[5317] <= 1'b1;
pika_color[5367] <= 1'b1;
pika_color[5421] <= 1'b1;
pika_color[5422] <= 1'b1;
pika_color[5431] <= 1'b1;
pika_color[5432] <= 1'b1;
pika_color[5482] <= 1'b1;
pika_color[5483] <= 1'b1;
pika_color[5537] <= 1'b1;
pika_color[5538] <= 1'b1;
pika_color[5546] <= 1'b1;
pika_color[5557] <= 1'b1;
pika_color[5558] <= 1'b1;
pika_color[5559] <= 1'b1;
pika_color[5598] <= 1'b1;
pika_color[5653] <= 1'b1;
pika_color[5654] <= 1'b1;
pika_color[5661] <= 1'b1;
pika_color[5671] <= 1'b1;
pika_color[5673] <= 1'b1;
pika_color[5674] <= 1'b1;
pika_color[5675] <= 1'b1;
pika_color[5698] <= 1'b1;
pika_color[5699] <= 1'b1;
pika_color[5713] <= 1'b1;
pika_color[5770] <= 1'b1;
pika_color[5776] <= 1'b1;
pika_color[5785] <= 1'b1;
pika_color[5789] <= 1'b1;
pika_color[5790] <= 1'b1;
pika_color[5791] <= 1'b1;
pika_color[5812] <= 1'b1;
pika_color[5814] <= 1'b1;
pika_color[5815] <= 1'b1;
pika_color[5816] <= 1'b1;
pika_color[5828] <= 1'b1;
pika_color[5885] <= 1'b1;
pika_color[5886] <= 1'b1;
pika_color[5891] <= 1'b1;
pika_color[5900] <= 1'b1;
pika_color[5904] <= 1'b1;
pika_color[5905] <= 1'b1;
pika_color[5906] <= 1'b1;
pika_color[5926] <= 1'b1;
pika_color[5930] <= 1'b1;
pika_color[5931] <= 1'b1;
pika_color[5932] <= 1'b1;
pika_color[5943] <= 1'b1;
pika_color[6002] <= 1'b1;
pika_color[6003] <= 1'b1;
pika_color[6006] <= 1'b1;
pika_color[6015] <= 1'b1;
pika_color[6016] <= 1'b1;
pika_color[6018] <= 1'b1;
pika_color[6019] <= 1'b1;
pika_color[6020] <= 1'b1;
pika_color[6021] <= 1'b1;
pika_color[6041] <= 1'b1;
pika_color[6046] <= 1'b1;
pika_color[6047] <= 1'b1;
pika_color[6058] <= 1'b1;
pika_color[6118] <= 1'b1;
pika_color[6119] <= 1'b1;
pika_color[6120] <= 1'b1;
pika_color[6121] <= 1'b1;
pika_color[6130] <= 1'b1;
pika_color[6131] <= 1'b1;
pika_color[6134] <= 1'b1;
pika_color[6136] <= 1'b1;
pika_color[6156] <= 1'b1;
pika_color[6157] <= 1'b1;
pika_color[6159] <= 1'b1;
pika_color[6160] <= 1'b1;
pika_color[6161] <= 1'b1;
pika_color[6162] <= 1'b1;
pika_color[6173] <= 1'b1;
pika_color[6234] <= 1'b1;
pika_color[6235] <= 1'b1;
pika_color[6246] <= 1'b1;
pika_color[6247] <= 1'b1;
pika_color[6249] <= 1'b1;
pika_color[6250] <= 1'b1;
pika_color[6271] <= 1'b1;
pika_color[6272] <= 1'b1;
pika_color[6274] <= 1'b1;
pika_color[6275] <= 1'b1;
pika_color[6276] <= 1'b1;
pika_color[6277] <= 1'b1;
pika_color[6288] <= 1'b1;
pika_color[6350] <= 1'b1;
pika_color[6362] <= 1'b1;
pika_color[6363] <= 1'b1;
pika_color[6364] <= 1'b1;
pika_color[6387] <= 1'b1;
pika_color[6388] <= 1'b1;
pika_color[6389] <= 1'b1;
pika_color[6390] <= 1'b1;
pika_color[6391] <= 1'b1;
pika_color[6403] <= 1'b1;
pika_color[6465] <= 1'b1;
pika_color[6503] <= 1'b1;
pika_color[6504] <= 1'b1;
pika_color[6505] <= 1'b1;
pika_color[6518] <= 1'b1;
pika_color[6580] <= 1'b1;
pika_color[6633] <= 1'b1;
pika_color[6695] <= 1'b1;
pika_color[6719] <= 1'b1;
pika_color[6720] <= 1'b1;
pika_color[6721] <= 1'b1;
pika_color[6722] <= 1'b1;
pika_color[6723] <= 1'b1;
pika_color[6748] <= 1'b1;
pika_color[6810] <= 1'b1;
pika_color[6835] <= 1'b1;
pika_color[6836] <= 1'b1;
pika_color[6837] <= 1'b1;
pika_color[6863] <= 1'b1;
pika_color[6925] <= 1'b1;
pika_color[6978] <= 1'b1;
pika_color[7040] <= 1'b1;
pika_color[7041] <= 1'b1;
pika_color[7093] <= 1'b1;
pika_color[7156] <= 1'b1;
pika_color[7208] <= 1'b1;
pika_color[7271] <= 1'b1;
pika_color[7272] <= 1'b1;
pika_color[7295] <= 1'b1;
pika_color[7296] <= 1'b1;
pika_color[7323] <= 1'b1;
pika_color[7386] <= 1'b1;
pika_color[7387] <= 1'b1;
pika_color[7409] <= 1'b1;
pika_color[7410] <= 1'b1;
pika_color[7412] <= 1'b1;
pika_color[7437] <= 1'b1;
pika_color[7438] <= 1'b1;
pika_color[7500] <= 1'b1;
pika_color[7501] <= 1'b1;
pika_color[7502] <= 1'b1;
pika_color[7503] <= 1'b1;
pika_color[7523] <= 1'b1;
pika_color[7524] <= 1'b1;
pika_color[7528] <= 1'b1;
pika_color[7552] <= 1'b1;
pika_color[7615] <= 1'b1;
pika_color[7618] <= 1'b1;
pika_color[7619] <= 1'b1;
pika_color[7638] <= 1'b1;
pika_color[7644] <= 1'b1;
pika_color[7666] <= 1'b1;
pika_color[7667] <= 1'b1;
pika_color[7728] <= 1'b1;
pika_color[7729] <= 1'b1;
pika_color[7730] <= 1'b1;
pika_color[7731] <= 1'b1;
pika_color[7732] <= 1'b1;
pika_color[7733] <= 1'b1;
pika_color[7734] <= 1'b1;
pika_color[7753] <= 1'b1;
pika_color[7759] <= 1'b1;
pika_color[7781] <= 1'b1;
pika_color[7842] <= 1'b1;
pika_color[7843] <= 1'b1;
pika_color[7849] <= 1'b1;
pika_color[7850] <= 1'b1;
pika_color[7851] <= 1'b1;
pika_color[7868] <= 1'b1;
pika_color[7870] <= 1'b1;
pika_color[7871] <= 1'b1;
pika_color[7872] <= 1'b1;
pika_color[7874] <= 1'b1;
pika_color[7896] <= 1'b1;
pika_color[7955] <= 1'b1;
pika_color[7956] <= 1'b1;
pika_color[7957] <= 1'b1;
pika_color[7966] <= 1'b1;
pika_color[7967] <= 1'b1;
pika_color[7983] <= 1'b1;
pika_color[7984] <= 1'b1;
pika_color[7988] <= 1'b1;
pika_color[7989] <= 1'b1;
pika_color[8011] <= 1'b1;
pika_color[8068] <= 1'b1;
pika_color[8069] <= 1'b1;
pika_color[8070] <= 1'b1;
pika_color[8082] <= 1'b1;
pika_color[8083] <= 1'b1;
pika_color[8098] <= 1'b1;
pika_color[8099] <= 1'b1;
pika_color[8103] <= 1'b1;
pika_color[8104] <= 1'b1;
pika_color[8125] <= 1'b1;
pika_color[8126] <= 1'b1;
pika_color[8183] <= 1'b1;
pika_color[8198] <= 1'b1;
pika_color[8199] <= 1'b1;
pika_color[8214] <= 1'b1;
pika_color[8215] <= 1'b1;
pika_color[8216] <= 1'b1;
pika_color[8217] <= 1'b1;
pika_color[8218] <= 1'b1;
pika_color[8239] <= 1'b1;
pika_color[8240] <= 1'b1;
pika_color[8241] <= 1'b1;
pika_color[8297] <= 1'b1;
pika_color[8314] <= 1'b1;
pika_color[8315] <= 1'b1;
pika_color[8353] <= 1'b1;
pika_color[8354] <= 1'b1;
pika_color[8356] <= 1'b1;
pika_color[8357] <= 1'b1;
pika_color[8412] <= 1'b1;
pika_color[8430] <= 1'b1;
pika_color[8431] <= 1'b1;
pika_color[8467] <= 1'b1;
pika_color[8468] <= 1'b1;
pika_color[8472] <= 1'b1;
pika_color[8473] <= 1'b1;
pika_color[8526] <= 1'b1;
pika_color[8546] <= 1'b1;
pika_color[8581] <= 1'b1;
pika_color[8582] <= 1'b1;
pika_color[8588] <= 1'b1;
pika_color[8641] <= 1'b1;
pika_color[8642] <= 1'b1;
pika_color[8662] <= 1'b1;
pika_color[8694] <= 1'b1;
pika_color[8695] <= 1'b1;
pika_color[8696] <= 1'b1;
pika_color[8703] <= 1'b1;
pika_color[8704] <= 1'b1;
pika_color[8757] <= 1'b1;
pika_color[8777] <= 1'b1;
pika_color[8778] <= 1'b1;
pika_color[8808] <= 1'b1;
pika_color[8809] <= 1'b1;
pika_color[8819] <= 1'b1;
pika_color[8872] <= 1'b1;
pika_color[8893] <= 1'b1;
pika_color[8894] <= 1'b1;
pika_color[8934] <= 1'b1;
pika_color[8935] <= 1'b1;
pika_color[8987] <= 1'b1;
pika_color[8988] <= 1'b1;
pika_color[9009] <= 1'b1;
pika_color[9050] <= 1'b1;
pika_color[9103] <= 1'b1;
pika_color[9104] <= 1'b1;
pika_color[9124] <= 1'b1;
pika_color[9125] <= 1'b1;
pika_color[9165] <= 1'b1;
pika_color[9219] <= 1'b1;
pika_color[9220] <= 1'b1;
pika_color[9240] <= 1'b1;
pika_color[9241] <= 1'b1;
pika_color[9280] <= 1'b1;
pika_color[9281] <= 1'b1;
pika_color[9335] <= 1'b1;
pika_color[9356] <= 1'b1;
pika_color[9357] <= 1'b1;
pika_color[9396] <= 1'b1;
pika_color[9451] <= 1'b1;
pika_color[9472] <= 1'b1;
pika_color[9473] <= 1'b1;
pika_color[9511] <= 1'b1;
pika_color[9566] <= 1'b1;
pika_color[9567] <= 1'b1;
pika_color[9588] <= 1'b1;
pika_color[9589] <= 1'b1;
pika_color[9608] <= 1'b1;
pika_color[9626] <= 1'b1;
pika_color[9682] <= 1'b1;
pika_color[9705] <= 1'b1;
pika_color[9723] <= 1'b1;
pika_color[9741] <= 1'b1;
pika_color[9797] <= 1'b1;
pika_color[9798] <= 1'b1;
pika_color[9838] <= 1'b1;
pika_color[9839] <= 1'b1;
pika_color[9856] <= 1'b1;
pika_color[9912] <= 1'b1;
pika_color[9913] <= 1'b1;
pika_color[9914] <= 1'b1;
pika_color[9954] <= 1'b1;
pika_color[9971] <= 1'b1;
pika_color[10027] <= 1'b1;
pika_color[10029] <= 1'b1;
pika_color[10030] <= 1'b1;
pika_color[10069] <= 1'b1;
pika_color[10070] <= 1'b1;
pika_color[10086] <= 1'b1;
pika_color[10142] <= 1'b1;
pika_color[10145] <= 1'b1;
pika_color[10146] <= 1'b1;
pika_color[10185] <= 1'b1;
pika_color[10201] <= 1'b1;
pika_color[10257] <= 1'b1;
pika_color[10261] <= 1'b1;
pika_color[10300] <= 1'b1;
pika_color[10316] <= 1'b1;
pika_color[10372] <= 1'b1;
pika_color[10376] <= 1'b1;
pika_color[10377] <= 1'b1;
pika_color[10415] <= 1'b1;
pika_color[10416] <= 1'b1;
pika_color[10431] <= 1'b1;
pika_color[10486] <= 1'b1;
pika_color[10487] <= 1'b1;
pika_color[10492] <= 1'b1;
pika_color[10531] <= 1'b1;
pika_color[10546] <= 1'b1;
pika_color[10601] <= 1'b1;
pika_color[10607] <= 1'b1;
pika_color[10608] <= 1'b1;
pika_color[10646] <= 1'b1;
pika_color[10647] <= 1'b1;
pika_color[10661] <= 1'b1;
pika_color[10716] <= 1'b1;
pika_color[10723] <= 1'b1;
pika_color[10762] <= 1'b1;
pika_color[10763] <= 1'b1;
pika_color[10776] <= 1'b1;
pika_color[10831] <= 1'b1;
pika_color[10878] <= 1'b1;
pika_color[10879] <= 1'b1;
pika_color[10880] <= 1'b1;
pika_color[10891] <= 1'b1;
pika_color[10945] <= 1'b1;
pika_color[10946] <= 1'b1;
pika_color[10995] <= 1'b1;
pika_color[11005] <= 1'b1;
pika_color[11006] <= 1'b1;
pika_color[11060] <= 1'b1;
pika_color[11110] <= 1'b1;
pika_color[11111] <= 1'b1;
pika_color[11112] <= 1'b1;
pika_color[11119] <= 1'b1;
pika_color[11120] <= 1'b1;
pika_color[11175] <= 1'b1;
pika_color[11227] <= 1'b1;
pika_color[11228] <= 1'b1;
pika_color[11233] <= 1'b1;
pika_color[11234] <= 1'b1;
pika_color[11290] <= 1'b1;
pika_color[11343] <= 1'b1;
pika_color[11344] <= 1'b1;
pika_color[11345] <= 1'b1;
pika_color[11346] <= 1'b1;
pika_color[11347] <= 1'b1;
pika_color[11348] <= 1'b1;
pika_color[11405] <= 1'b1;
pika_color[11461] <= 1'b1;
pika_color[11520] <= 1'b1;
pika_color[11576] <= 1'b1;
pika_color[11577] <= 1'b1;
pika_color[11635] <= 1'b1;
pika_color[11692] <= 1'b1;
pika_color[11750] <= 1'b1;
pika_color[11807] <= 1'b1;
pika_color[11865] <= 1'b1;
pika_color[11922] <= 1'b1;
pika_color[11980] <= 1'b1;
pika_color[12037] <= 1'b1;
pika_color[12095] <= 1'b1;
pika_color[12152] <= 1'b1;
pika_color[12210] <= 1'b1;
pika_color[12267] <= 1'b1;
pika_color[12325] <= 1'b1;
pika_color[12382] <= 1'b1;
pika_color[12440] <= 1'b1;
pika_color[12497] <= 1'b1;
pika_color[12555] <= 1'b1;
pika_color[12612] <= 1'b1;
pika_color[12670] <= 1'b1;
pika_color[12671] <= 1'b1;
pika_color[12727] <= 1'b1;
pika_color[12786] <= 1'b1;
pika_color[12842] <= 1'b1;
pika_color[12901] <= 1'b1;
pika_color[12957] <= 1'b1;
pika_color[13016] <= 1'b1;
pika_color[13072] <= 1'b1;
pika_color[13131] <= 1'b1;
pika_color[13187] <= 1'b1;
pika_color[13246] <= 1'b1;
pika_color[13302] <= 1'b1;
pika_color[13361] <= 1'b1;
pika_color[13362] <= 1'b1;
pika_color[13417] <= 1'b1;
pika_color[13477] <= 1'b1;
pika_color[13532] <= 1'b1;
pika_color[13592] <= 1'b1;
pika_color[13593] <= 1'b1;
pika_color[13647] <= 1'b1;
pika_color[13708] <= 1'b1;
pika_color[13762] <= 1'b1;
pika_color[13823] <= 1'b1;
pika_color[13877] <= 1'b1;
pika_color[13938] <= 1'b1;
pika_color[13939] <= 1'b1;
pika_color[13991] <= 1'b1;
pika_color[13992] <= 1'b1;
pika_color[14054] <= 1'b1;
pika_color[14106] <= 1'b1;
pika_color[14169] <= 1'b1;
pika_color[14170] <= 1'b1;
pika_color[14220] <= 1'b1;
pika_color[14221] <= 1'b1;
pika_color[14285] <= 1'b1;
pika_color[14334] <= 1'b1;
pika_color[14335] <= 1'b1;
pika_color[14400] <= 1'b1;
pika_color[14401] <= 1'b1;
pika_color[14448] <= 1'b1;
pika_color[14449] <= 1'b1;
pika_color[14516] <= 1'b1;
pika_color[14517] <= 1'b1;
pika_color[14518] <= 1'b1;
pika_color[14519] <= 1'b1;
pika_color[14532] <= 1'b1;
pika_color[14533] <= 1'b1;
pika_color[14534] <= 1'b1;
pika_color[14535] <= 1'b1;
pika_color[14536] <= 1'b1;
pika_color[14537] <= 1'b1;
pika_color[14538] <= 1'b1;
pika_color[14539] <= 1'b1;
pika_color[14540] <= 1'b1;
pika_color[14541] <= 1'b1;
pika_color[14542] <= 1'b1;
pika_color[14543] <= 1'b1;
pika_color[14544] <= 1'b1;
pika_color[14545] <= 1'b1;
pika_color[14546] <= 1'b1;
pika_color[14562] <= 1'b1;
pika_color[14563] <= 1'b1;
pika_color[14634] <= 1'b1;
pika_color[14635] <= 1'b1;
pika_color[14636] <= 1'b1;
pika_color[14637] <= 1'b1;
pika_color[14647] <= 1'b1;
pika_color[14661] <= 1'b1;
pika_color[14662] <= 1'b1;
pika_color[14663] <= 1'b1;
pika_color[14664] <= 1'b1;
pika_color[14665] <= 1'b1;
pika_color[14676] <= 1'b1;
pika_color[14677] <= 1'b1;
pika_color[14751] <= 1'b1;
pika_color[14761] <= 1'b1;
pika_color[14762] <= 1'b1;
pika_color[14780] <= 1'b1;
pika_color[14790] <= 1'b1;
pika_color[14791] <= 1'b1;
pika_color[14866] <= 1'b1;
pika_color[14876] <= 1'b1;
pika_color[14895] <= 1'b1;
pika_color[14896] <= 1'b1;
pika_color[14905] <= 1'b1;
pika_color[14981] <= 1'b1;
pika_color[14982] <= 1'b1;
pika_color[14990] <= 1'b1;
pika_color[14991] <= 1'b1;
pika_color[15011] <= 1'b1;
pika_color[15020] <= 1'b1;
pika_color[15097] <= 1'b1;
pika_color[15098] <= 1'b1;
pika_color[15099] <= 1'b1;
pika_color[15100] <= 1'b1;
pika_color[15101] <= 1'b1;
pika_color[15102] <= 1'b1;
pika_color[15103] <= 1'b1;
pika_color[15104] <= 1'b1;
pika_color[15126] <= 1'b1;
pika_color[15127] <= 1'b1;
pika_color[15135] <= 1'b1;
pika_color[15242] <= 1'b1;
pika_color[15243] <= 1'b1;
pika_color[15244] <= 1'b1;
pika_color[15250] <= 1'b1;
pika_color[15251] <= 1'b1;
pika_color[15359] <= 1'b1;
pika_color[15360] <= 1'b1;
pika_color[15366] <= 1'b1;
pika_color[15367] <= 1'b1;
pika_color[15475] <= 1'b1;
pika_color[15476] <= 1'b1;
pika_color[15482] <= 1'b1;
pika_color[15483] <= 1'b1;
pika_color[15591] <= 1'b1;
pika_color[15598] <= 1'b1;
pika_color[15599] <= 1'b1;
pika_color[15706] <= 1'b1;
pika_color[15714] <= 1'b1;
pika_color[15715] <= 1'b1;
pika_color[15821] <= 1'b1;
pika_color[15831] <= 1'b1;
pika_color[15936] <= 1'b1;
pika_color[15946] <= 1'b1;
pika_color[16051] <= 1'b1;
pika_color[16052] <= 1'b1;
pika_color[16061] <= 1'b1;
pika_color[16167] <= 1'b1;
pika_color[16168] <= 1'b1;
pika_color[16169] <= 1'b1;
pika_color[16170] <= 1'b1;
pika_color[16174] <= 1'b1;
pika_color[16175] <= 1'b1;
pika_color[16176] <= 1'b1;
pika_color[16285] <= 1'b1;
pika_color[16286] <= 1'b1;
pika_color[16287] <= 1'b1;
pika_color[16288] <= 1'b1;
pika_color[16289] <= 1'b1;

end
		default:;
	endcase
	end
	
	
endmodule