module left_Score(input Reset, frame_clk, output [1374:0] score_bar_left);
	always_comb
	 begin
	score_bar_left[279] <= 1'b1;
score_bar_left[280] <= 1'b1;
score_bar_left[281] <= 1'b1;
score_bar_left[282] <= 1'b1;
score_bar_left[283] <= 1'b1;
score_bar_left[284] <= 1'b1;
score_bar_left[333] <= 1'b1;
score_bar_left[334] <= 1'b1;
score_bar_left[335] <= 1'b1;
score_bar_left[338] <= 1'b1;
score_bar_left[339] <= 1'b1;
score_bar_left[387] <= 1'b1;
score_bar_left[388] <= 1'b1;
score_bar_left[442] <= 1'b1;
score_bar_left[443] <= 1'b1;
score_bar_left[497] <= 1'b1;
score_bar_left[498] <= 1'b1;
score_bar_left[510] <= 1'b1;
score_bar_left[511] <= 1'b1;
score_bar_left[512] <= 1'b1;
score_bar_left[513] <= 1'b1;
score_bar_left[514] <= 1'b1;
score_bar_left[519] <= 1'b1;
score_bar_left[520] <= 1'b1;
score_bar_left[521] <= 1'b1;
score_bar_left[522] <= 1'b1;
score_bar_left[523] <= 1'b1;
score_bar_left[529] <= 1'b1;
score_bar_left[531] <= 1'b1;
score_bar_left[532] <= 1'b1;
score_bar_left[533] <= 1'b1;
score_bar_left[538] <= 1'b1;
score_bar_left[539] <= 1'b1;
score_bar_left[540] <= 1'b1;
score_bar_left[541] <= 1'b1;
score_bar_left[546] <= 1'b1;
score_bar_left[547] <= 1'b1;
score_bar_left[553] <= 1'b1;
score_bar_left[554] <= 1'b1;
score_bar_left[564] <= 1'b1;
score_bar_left[565] <= 1'b1;
score_bar_left[569] <= 1'b1;
score_bar_left[573] <= 1'b1;
score_bar_left[574] <= 1'b1;
score_bar_left[578] <= 1'b1;
score_bar_left[579] <= 1'b1;
score_bar_left[584] <= 1'b1;
score_bar_left[585] <= 1'b1;
score_bar_left[586] <= 1'b1;
score_bar_left[592] <= 1'b1;
score_bar_left[593] <= 1'b1;
score_bar_left[596] <= 1'b1;
score_bar_left[597] <= 1'b1;
score_bar_left[601] <= 1'b1;
score_bar_left[602] <= 1'b1;
score_bar_left[609] <= 1'b1;
score_bar_left[610] <= 1'b1;
score_bar_left[611] <= 1'b1;
score_bar_left[618] <= 1'b1;
score_bar_left[619] <= 1'b1;
score_bar_left[627] <= 1'b1;
score_bar_left[628] <= 1'b1;
score_bar_left[634] <= 1'b1;
score_bar_left[635] <= 1'b1;
score_bar_left[639] <= 1'b1;
score_bar_left[640] <= 1'b1;
score_bar_left[646] <= 1'b1;
score_bar_left[647] <= 1'b1;
score_bar_left[652] <= 1'b1;
score_bar_left[653] <= 1'b1;
score_bar_left[666] <= 1'b1;
score_bar_left[667] <= 1'b1;
score_bar_left[668] <= 1'b1;
score_bar_left[673] <= 1'b1;
score_bar_left[682] <= 1'b1;
score_bar_left[690] <= 1'b1;
score_bar_left[694] <= 1'b1;
score_bar_left[700] <= 1'b1;
score_bar_left[701] <= 1'b1;
score_bar_left[708] <= 1'b1;
score_bar_left[709] <= 1'b1;
score_bar_left[723] <= 1'b1;
score_bar_left[724] <= 1'b1;
score_bar_left[727] <= 1'b1;
score_bar_left[728] <= 1'b1;
score_bar_left[736] <= 1'b1;
score_bar_left[737] <= 1'b1;
score_bar_left[745] <= 1'b1;
score_bar_left[746] <= 1'b1;
score_bar_left[749] <= 1'b1;
score_bar_left[755] <= 1'b1;
score_bar_left[756] <= 1'b1;
score_bar_left[757] <= 1'b1;
score_bar_left[758] <= 1'b1;
score_bar_left[759] <= 1'b1;
score_bar_left[760] <= 1'b1;
score_bar_left[761] <= 1'b1;
score_bar_left[762] <= 1'b1;
score_bar_left[763] <= 1'b1;
score_bar_left[764] <= 1'b1;
score_bar_left[779] <= 1'b1;
score_bar_left[780] <= 1'b1;
score_bar_left[782] <= 1'b1;
score_bar_left[783] <= 1'b1;
score_bar_left[791] <= 1'b1;
score_bar_left[792] <= 1'b1;
score_bar_left[800] <= 1'b1;
score_bar_left[801] <= 1'b1;
score_bar_left[804] <= 1'b1;
score_bar_left[810] <= 1'b1;
score_bar_left[811] <= 1'b1;
score_bar_left[834] <= 1'b1;
score_bar_left[835] <= 1'b1;
score_bar_left[838] <= 1'b1;
score_bar_left[847] <= 1'b1;
score_bar_left[855] <= 1'b1;
score_bar_left[859] <= 1'b1;
score_bar_left[865] <= 1'b1;
score_bar_left[866] <= 1'b1;
score_bar_left[882] <= 1'b1;
score_bar_left[889] <= 1'b1;
score_bar_left[890] <= 1'b1;
score_bar_left[893] <= 1'b1;
score_bar_left[894] <= 1'b1;
score_bar_left[902] <= 1'b1;
score_bar_left[903] <= 1'b1;
score_bar_left[909] <= 1'b1;
score_bar_left[910] <= 1'b1;
score_bar_left[914] <= 1'b1;
score_bar_left[921] <= 1'b1;
score_bar_left[922] <= 1'b1;
score_bar_left[937] <= 1'b1;
score_bar_left[938] <= 1'b1;
score_bar_left[942] <= 1'b1;
score_bar_left[943] <= 1'b1;
score_bar_left[944] <= 1'b1;
score_bar_left[949] <= 1'b1;
score_bar_left[950] <= 1'b1;
score_bar_left[954] <= 1'b1;
score_bar_left[958] <= 1'b1;
score_bar_left[959] <= 1'b1;
score_bar_left[963] <= 1'b1;
score_bar_left[964] <= 1'b1;
score_bar_left[969] <= 1'b1;
score_bar_left[977] <= 1'b1;
score_bar_left[978] <= 1'b1;
score_bar_left[982] <= 1'b1;
score_bar_left[983] <= 1'b1;
score_bar_left[986] <= 1'b1;
score_bar_left[987] <= 1'b1;
score_bar_left[993] <= 1'b1;
score_bar_left[994] <= 1'b1;
score_bar_left[995] <= 1'b1;
score_bar_left[996] <= 1'b1;
score_bar_left[997] <= 1'b1;
score_bar_left[1005] <= 1'b1;
score_bar_left[1006] <= 1'b1;
score_bar_left[1007] <= 1'b1;
score_bar_left[1008] <= 1'b1;
score_bar_left[1009] <= 1'b1;
score_bar_left[1014] <= 1'b1;
score_bar_left[1015] <= 1'b1;
score_bar_left[1016] <= 1'b1;
score_bar_left[1017] <= 1'b1;
score_bar_left[1018] <= 1'b1;
score_bar_left[1024] <= 1'b1;
score_bar_left[1033] <= 1'b1;
score_bar_left[1034] <= 1'b1;
score_bar_left[1035] <= 1'b1;
score_bar_left[1036] <= 1'b1;
score_bar_left[1037] <= 1'b1;
score_bar_left[1041] <= 1'b1;
score_bar_left[1042] <= 1'b1;


	 end
endmodule