module start_screen_text_display(input Reset, frame_clk, 
														input logic [7:0] keycode,
														output [20999:0] startscreen);
														
								
	 enum logic [3:0] {Halted, Normal} State, Next_state;
	 logic display_text;
	 always_ff @ (posedge frame_clk )
    begin
		if(Reset)
			State <= Halted;
		else
			State <= Next_state;
    end
	 
	 always_comb
	 begin
		Next_state = State;
		display_text = 1'b1;
		unique case(State)
			Halted:
			begin
				display_text = 1'b1;
				if(keycode == 8'h2c)
					Next_state = Normal;
			end
			Normal:
				display_text = 1'b0;
		endcase
					
	 end
	 
	 always_comb
	 begin
	 startscreen <= 1'b0;
	 if(display_text == 1'b1)
	 begin
		startscreen[2527] <= 1'b1;
startscreen[2528] <= 1'b1;
startscreen[2529] <= 1'b1;
startscreen[2530] <= 1'b1;
startscreen[2531] <= 1'b1;
startscreen[2532] <= 1'b1;
startscreen[2533] <= 1'b1;
startscreen[2534] <= 1'b1;
startscreen[2535] <= 1'b1;
startscreen[2536] <= 1'b1;
startscreen[2537] <= 1'b1;
startscreen[2538] <= 1'b1;
startscreen[2539] <= 1'b1;
startscreen[2540] <= 1'b1;
startscreen[2656] <= 1'b1;
startscreen[2657] <= 1'b1;
startscreen[2658] <= 1'b1;
startscreen[2659] <= 1'b1;
startscreen[2660] <= 1'b1;
startscreen[2661] <= 1'b1;
startscreen[2662] <= 1'b1;
startscreen[2663] <= 1'b1;
startscreen[2852] <= 1'b1;
startscreen[2853] <= 1'b1;
startscreen[2854] <= 1'b1;
startscreen[2855] <= 1'b1;
startscreen[2856] <= 1'b1;
startscreen[2857] <= 1'b1;
startscreen[2858] <= 1'b1;
startscreen[2859] <= 1'b1;
startscreen[2947] <= 1'b1;
startscreen[2949] <= 1'b1;
startscreen[2950] <= 1'b1;
startscreen[2951] <= 1'b1;
startscreen[2952] <= 1'b1;
startscreen[2953] <= 1'b1;
startscreen[2954] <= 1'b1;
startscreen[2955] <= 1'b1;
startscreen[2956] <= 1'b1;
startscreen[2957] <= 1'b1;
startscreen[2958] <= 1'b1;
startscreen[2959] <= 1'b1;
startscreen[2960] <= 1'b1;
startscreen[2961] <= 1'b1;
startscreen[2962] <= 1'b1;
startscreen[3073] <= 1'b1;
startscreen[3076] <= 1'b1;
startscreen[3077] <= 1'b1;
startscreen[3078] <= 1'b1;
startscreen[3079] <= 1'b1;
startscreen[3080] <= 1'b1;
startscreen[3081] <= 1'b1;
startscreen[3082] <= 1'b1;
startscreen[3083] <= 1'b1;
startscreen[3084] <= 1'b1;
startscreen[3085] <= 1'b1;
startscreen[3086] <= 1'b1;
startscreen[3269] <= 1'b1;
startscreen[3270] <= 1'b1;
startscreen[3271] <= 1'b1;
startscreen[3273] <= 1'b1;
startscreen[3274] <= 1'b1;
startscreen[3275] <= 1'b1;
startscreen[3278] <= 1'b1;
startscreen[3279] <= 1'b1;
startscreen[3280] <= 1'b1;
startscreen[3281] <= 1'b1;
startscreen[3282] <= 1'b1;
startscreen[3367] <= 1'b1;
startscreen[3368] <= 1'b1;
startscreen[3369] <= 1'b1;
startscreen[3371] <= 1'b1;
startscreen[3372] <= 1'b1;
startscreen[3373] <= 1'b1;
startscreen[3375] <= 1'b1;
startscreen[3376] <= 1'b1;
startscreen[3381] <= 1'b1;
startscreen[3382] <= 1'b1;
startscreen[3383] <= 1'b1;
startscreen[3491] <= 1'b1;
startscreen[3492] <= 1'b1;
startscreen[3494] <= 1'b1;
startscreen[3495] <= 1'b1;
startscreen[3498] <= 1'b1;
startscreen[3500] <= 1'b1;
startscreen[3501] <= 1'b1;
startscreen[3502] <= 1'b1;
startscreen[3503] <= 1'b1;
startscreen[3504] <= 1'b1;
startscreen[3505] <= 1'b1;
startscreen[3506] <= 1'b1;
startscreen[3631] <= 1'b1;
startscreen[3632] <= 1'b1;
startscreen[3687] <= 1'b1;
startscreen[3688] <= 1'b1;
startscreen[3689] <= 1'b1;
startscreen[3690] <= 1'b1;
startscreen[3691] <= 1'b1;
startscreen[3692] <= 1'b1;
startscreen[3693] <= 1'b1;
startscreen[3694] <= 1'b1;
startscreen[3695] <= 1'b1;
startscreen[3696] <= 1'b1;
startscreen[3697] <= 1'b1;
startscreen[3698] <= 1'b1;
startscreen[3699] <= 1'b1;
startscreen[3701] <= 1'b1;
startscreen[3702] <= 1'b1;
startscreen[3712] <= 1'b1;
startscreen[3713] <= 1'b1;
startscreen[3769] <= 1'b1;
startscreen[3770] <= 1'b1;
startscreen[3787] <= 1'b1;
startscreen[3788] <= 1'b1;
startscreen[3790] <= 1'b1;
startscreen[3791] <= 1'b1;
startscreen[3792] <= 1'b1;
startscreen[3793] <= 1'b1;
startscreen[3794] <= 1'b1;
startscreen[3795] <= 1'b1;
startscreen[3796] <= 1'b1;
startscreen[3797] <= 1'b1;
startscreen[3798] <= 1'b1;
startscreen[3799] <= 1'b1;
startscreen[3800] <= 1'b1;
startscreen[3801] <= 1'b1;
startscreen[3804] <= 1'b1;
startscreen[3910] <= 1'b1;
startscreen[3911] <= 1'b1;
startscreen[3912] <= 1'b1;
startscreen[3913] <= 1'b1;
startscreen[3914] <= 1'b1;
startscreen[3915] <= 1'b1;
startscreen[3916] <= 1'b1;
startscreen[3917] <= 1'b1;
startscreen[3921] <= 1'b1;
startscreen[3922] <= 1'b1;
startscreen[3923] <= 1'b1;
startscreen[3924] <= 1'b1;
startscreen[3925] <= 1'b1;
startscreen[3926] <= 1'b1;
startscreen[4049] <= 1'b1;
startscreen[4050] <= 1'b1;
startscreen[4051] <= 1'b1;
startscreen[4052] <= 1'b1;
startscreen[4106] <= 1'b1;
startscreen[4107] <= 1'b1;
startscreen[4109] <= 1'b1;
startscreen[4110] <= 1'b1;
startscreen[4111] <= 1'b1;
startscreen[4112] <= 1'b1;
startscreen[4113] <= 1'b1;
startscreen[4117] <= 1'b1;
startscreen[4118] <= 1'b1;
startscreen[4119] <= 1'b1;
startscreen[4120] <= 1'b1;
startscreen[4121] <= 1'b1;
startscreen[4122] <= 1'b1;
startscreen[4130] <= 1'b1;
startscreen[4131] <= 1'b1;
startscreen[4133] <= 1'b1;
startscreen[4187] <= 1'b1;
startscreen[4188] <= 1'b1;
startscreen[4189] <= 1'b1;
startscreen[4190] <= 1'b1;
startscreen[4207] <= 1'b1;
startscreen[4208] <= 1'b1;
startscreen[4209] <= 1'b1;
startscreen[4210] <= 1'b1;
startscreen[4223] <= 1'b1;
startscreen[4224] <= 1'b1;
startscreen[4225] <= 1'b1;
startscreen[4329] <= 1'b1;
startscreen[4330] <= 1'b1;
startscreen[4332] <= 1'b1;
startscreen[4333] <= 1'b1;
startscreen[4334] <= 1'b1;
startscreen[4344] <= 1'b1;
startscreen[4345] <= 1'b1;
startscreen[4346] <= 1'b1;
startscreen[4469] <= 1'b1;
startscreen[4471] <= 1'b1;
startscreen[4472] <= 1'b1;
startscreen[4525] <= 1'b1;
startscreen[4526] <= 1'b1;
startscreen[4527] <= 1'b1;
startscreen[4528] <= 1'b1;
startscreen[4529] <= 1'b1;
startscreen[4540] <= 1'b1;
startscreen[4541] <= 1'b1;
startscreen[4542] <= 1'b1;
startscreen[4550] <= 1'b1;
startscreen[4551] <= 1'b1;
startscreen[4552] <= 1'b1;
startscreen[4553] <= 1'b1;
startscreen[4607] <= 1'b1;
startscreen[4608] <= 1'b1;
startscreen[4610] <= 1'b1;
startscreen[4627] <= 1'b1;
startscreen[4628] <= 1'b1;
startscreen[4629] <= 1'b1;
startscreen[4630] <= 1'b1;
startscreen[4642] <= 1'b1;
startscreen[4643] <= 1'b1;
startscreen[4752] <= 1'b1;
startscreen[4765] <= 1'b1;
startscreen[4766] <= 1'b1;
startscreen[4889] <= 1'b1;
startscreen[4891] <= 1'b1;
startscreen[4892] <= 1'b1;
startscreen[4944] <= 1'b1;
startscreen[4945] <= 1'b1;
startscreen[4946] <= 1'b1;
startscreen[4947] <= 1'b1;
startscreen[4948] <= 1'b1;
startscreen[4970] <= 1'b1;
startscreen[4972] <= 1'b1;
startscreen[4973] <= 1'b1;
startscreen[5027] <= 1'b1;
startscreen[5028] <= 1'b1;
startscreen[5029] <= 1'b1;
startscreen[5030] <= 1'b1;
startscreen[5047] <= 1'b1;
startscreen[5048] <= 1'b1;
startscreen[5050] <= 1'b1;
startscreen[5063] <= 1'b1;
startscreen[5065] <= 1'b1;
startscreen[5066] <= 1'b1;
startscreen[5168] <= 1'b1;
startscreen[5170] <= 1'b1;
startscreen[5171] <= 1'b1;
startscreen[5309] <= 1'b1;
startscreen[5310] <= 1'b1;
startscreen[5311] <= 1'b1;
startscreen[5312] <= 1'b1;
startscreen[5364] <= 1'b1;
startscreen[5366] <= 1'b1;
startscreen[5367] <= 1'b1;
startscreen[5390] <= 1'b1;
startscreen[5393] <= 1'b1;
startscreen[5447] <= 1'b1;
startscreen[5448] <= 1'b1;
startscreen[5450] <= 1'b1;
startscreen[5467] <= 1'b1;
startscreen[5468] <= 1'b1;
startscreen[5469] <= 1'b1;
startscreen[5470] <= 1'b1;
startscreen[5483] <= 1'b1;
startscreen[5484] <= 1'b1;
startscreen[5485] <= 1'b1;
startscreen[5486] <= 1'b1;
startscreen[5588] <= 1'b1;
startscreen[5591] <= 1'b1;
startscreen[5730] <= 1'b1;
startscreen[5731] <= 1'b1;
startscreen[5732] <= 1'b1;
startscreen[5784] <= 1'b1;
startscreen[5786] <= 1'b1;
startscreen[5787] <= 1'b1;
startscreen[5810] <= 1'b1;
startscreen[5811] <= 1'b1;
startscreen[5812] <= 1'b1;
startscreen[5813] <= 1'b1;
startscreen[5867] <= 1'b1;
startscreen[5868] <= 1'b1;
startscreen[5870] <= 1'b1;
startscreen[5887] <= 1'b1;
startscreen[5888] <= 1'b1;
startscreen[5890] <= 1'b1;
startscreen[5904] <= 1'b1;
startscreen[5905] <= 1'b1;
startscreen[5906] <= 1'b1;
startscreen[6008] <= 1'b1;
startscreen[6009] <= 1'b1;
startscreen[6010] <= 1'b1;
startscreen[6011] <= 1'b1;
startscreen[6150] <= 1'b1;
startscreen[6152] <= 1'b1;
startscreen[6204] <= 1'b1;
startscreen[6206] <= 1'b1;
startscreen[6207] <= 1'b1;
startscreen[6230] <= 1'b1;
startscreen[6233] <= 1'b1;
startscreen[6287] <= 1'b1;
startscreen[6289] <= 1'b1;
startscreen[6290] <= 1'b1;
startscreen[6307] <= 1'b1;
startscreen[6308] <= 1'b1;
startscreen[6309] <= 1'b1;
startscreen[6310] <= 1'b1;
startscreen[6324] <= 1'b1;
startscreen[6325] <= 1'b1;
startscreen[6326] <= 1'b1;
startscreen[6333] <= 1'b1;
startscreen[6334] <= 1'b1;
startscreen[6335] <= 1'b1;
startscreen[6336] <= 1'b1;
startscreen[6342] <= 1'b1;
startscreen[6343] <= 1'b1;
startscreen[6344] <= 1'b1;
startscreen[6355] <= 1'b1;
startscreen[6356] <= 1'b1;
startscreen[6357] <= 1'b1;
startscreen[6358] <= 1'b1;
startscreen[6359] <= 1'b1;
startscreen[6360] <= 1'b1;
startscreen[6361] <= 1'b1;
startscreen[6362] <= 1'b1;
startscreen[6379] <= 1'b1;
startscreen[6380] <= 1'b1;
startscreen[6381] <= 1'b1;
startscreen[6382] <= 1'b1;
startscreen[6383] <= 1'b1;
startscreen[6384] <= 1'b1;
startscreen[6385] <= 1'b1;
startscreen[6400] <= 1'b1;
startscreen[6401] <= 1'b1;
startscreen[6402] <= 1'b1;
startscreen[6403] <= 1'b1;
startscreen[6404] <= 1'b1;
startscreen[6405] <= 1'b1;
startscreen[6428] <= 1'b1;
startscreen[6430] <= 1'b1;
startscreen[6431] <= 1'b1;
startscreen[6454] <= 1'b1;
startscreen[6455] <= 1'b1;
startscreen[6456] <= 1'b1;
startscreen[6457] <= 1'b1;
startscreen[6463] <= 1'b1;
startscreen[6464] <= 1'b1;
startscreen[6465] <= 1'b1;
startscreen[6466] <= 1'b1;
startscreen[6467] <= 1'b1;
startscreen[6468] <= 1'b1;
startscreen[6469] <= 1'b1;
startscreen[6488] <= 1'b1;
startscreen[6489] <= 1'b1;
startscreen[6490] <= 1'b1;
startscreen[6491] <= 1'b1;
startscreen[6492] <= 1'b1;
startscreen[6493] <= 1'b1;
startscreen[6494] <= 1'b1;
startscreen[6514] <= 1'b1;
startscreen[6515] <= 1'b1;
startscreen[6516] <= 1'b1;
startscreen[6517] <= 1'b1;
startscreen[6518] <= 1'b1;
startscreen[6519] <= 1'b1;
startscreen[6520] <= 1'b1;
startscreen[6521] <= 1'b1;
startscreen[6534] <= 1'b1;
startscreen[6535] <= 1'b1;
startscreen[6536] <= 1'b1;
startscreen[6537] <= 1'b1;
startscreen[6538] <= 1'b1;
startscreen[6539] <= 1'b1;
startscreen[6540] <= 1'b1;
startscreen[6541] <= 1'b1;
startscreen[6542] <= 1'b1;
startscreen[6564] <= 1'b1;
startscreen[6565] <= 1'b1;
startscreen[6566] <= 1'b1;
startscreen[6567] <= 1'b1;
startscreen[6568] <= 1'b1;
startscreen[6570] <= 1'b1;
startscreen[6572] <= 1'b1;
startscreen[6573] <= 1'b1;
startscreen[6575] <= 1'b1;
startscreen[6577] <= 1'b1;
startscreen[6578] <= 1'b1;
startscreen[6590] <= 1'b1;
startscreen[6591] <= 1'b1;
startscreen[6592] <= 1'b1;
startscreen[6593] <= 1'b1;
startscreen[6594] <= 1'b1;
startscreen[6595] <= 1'b1;
startscreen[6596] <= 1'b1;
startscreen[6597] <= 1'b1;
startscreen[6624] <= 1'b1;
startscreen[6626] <= 1'b1;
startscreen[6627] <= 1'b1;
startscreen[6646] <= 1'b1;
startscreen[6648] <= 1'b1;
startscreen[6650] <= 1'b1;
startscreen[6653] <= 1'b1;
startscreen[6654] <= 1'b1;
startscreen[6656] <= 1'b1;
startscreen[6657] <= 1'b1;
startscreen[6670] <= 1'b1;
startscreen[6671] <= 1'b1;
startscreen[6672] <= 1'b1;
startscreen[6673] <= 1'b1;
startscreen[6674] <= 1'b1;
startscreen[6675] <= 1'b1;
startscreen[6676] <= 1'b1;
startscreen[6677] <= 1'b1;
startscreen[6690] <= 1'b1;
startscreen[6692] <= 1'b1;
startscreen[6693] <= 1'b1;
startscreen[6698] <= 1'b1;
startscreen[6699] <= 1'b1;
startscreen[6700] <= 1'b1;
startscreen[6701] <= 1'b1;
startscreen[6703] <= 1'b1;
startscreen[6704] <= 1'b1;
startscreen[6705] <= 1'b1;
startscreen[6706] <= 1'b1;
startscreen[6707] <= 1'b1;
startscreen[6708] <= 1'b1;
startscreen[6709] <= 1'b1;
startscreen[6711] <= 1'b1;
startscreen[6712] <= 1'b1;
startscreen[6713] <= 1'b1;
startscreen[6715] <= 1'b1;
startscreen[6716] <= 1'b1;
startscreen[6717] <= 1'b1;
startscreen[6727] <= 1'b1;
startscreen[6728] <= 1'b1;
startscreen[6729] <= 1'b1;
startscreen[6730] <= 1'b1;
startscreen[6744] <= 1'b1;
startscreen[6745] <= 1'b1;
startscreen[6746] <= 1'b1;
startscreen[6753] <= 1'b1;
startscreen[6754] <= 1'b1;
startscreen[6755] <= 1'b1;
startscreen[6756] <= 1'b1;
startscreen[6760] <= 1'b1;
startscreen[6762] <= 1'b1;
startscreen[6763] <= 1'b1;
startscreen[6765] <= 1'b1;
startscreen[6773] <= 1'b1;
startscreen[6774] <= 1'b1;
startscreen[6776] <= 1'b1;
startscreen[6777] <= 1'b1;
startscreen[6780] <= 1'b1;
startscreen[6781] <= 1'b1;
startscreen[6782] <= 1'b1;
startscreen[6783] <= 1'b1;
startscreen[6784] <= 1'b1;
startscreen[6797] <= 1'b1;
startscreen[6799] <= 1'b1;
startscreen[6800] <= 1'b1;
startscreen[6801] <= 1'b1;
startscreen[6802] <= 1'b1;
startscreen[6803] <= 1'b1;
startscreen[6804] <= 1'b1;
startscreen[6805] <= 1'b1;
startscreen[6807] <= 1'b1;
startscreen[6820] <= 1'b1;
startscreen[6821] <= 1'b1;
startscreen[6823] <= 1'b1;
startscreen[6824] <= 1'b1;
startscreen[6825] <= 1'b1;
startscreen[6826] <= 1'b1;
startscreen[6827] <= 1'b1;
startscreen[6828] <= 1'b1;
startscreen[6848] <= 1'b1;
startscreen[6850] <= 1'b1;
startscreen[6851] <= 1'b1;
startscreen[6874] <= 1'b1;
startscreen[6875] <= 1'b1;
startscreen[6877] <= 1'b1;
startscreen[6881] <= 1'b1;
startscreen[6882] <= 1'b1;
startscreen[6885] <= 1'b1;
startscreen[6886] <= 1'b1;
startscreen[6889] <= 1'b1;
startscreen[6891] <= 1'b1;
startscreen[6905] <= 1'b1;
startscreen[6907] <= 1'b1;
startscreen[6908] <= 1'b1;
startscreen[6910] <= 1'b1;
startscreen[6911] <= 1'b1;
startscreen[6912] <= 1'b1;
startscreen[6913] <= 1'b1;
startscreen[6914] <= 1'b1;
startscreen[6915] <= 1'b1;
startscreen[6916] <= 1'b1;
startscreen[6932] <= 1'b1;
startscreen[6933] <= 1'b1;
startscreen[6934] <= 1'b1;
startscreen[6935] <= 1'b1;
startscreen[6936] <= 1'b1;
startscreen[6937] <= 1'b1;
startscreen[6938] <= 1'b1;
startscreen[6939] <= 1'b1;
startscreen[6940] <= 1'b1;
startscreen[6941] <= 1'b1;
startscreen[6942] <= 1'b1;
startscreen[6943] <= 1'b1;
startscreen[6952] <= 1'b1;
startscreen[6953] <= 1'b1;
startscreen[6954] <= 1'b1;
startscreen[6956] <= 1'b1;
startscreen[6957] <= 1'b1;
startscreen[6958] <= 1'b1;
startscreen[6959] <= 1'b1;
startscreen[6960] <= 1'b1;
startscreen[6962] <= 1'b1;
startscreen[6963] <= 1'b1;
startscreen[6964] <= 1'b1;
startscreen[6984] <= 1'b1;
startscreen[6987] <= 1'b1;
startscreen[6989] <= 1'b1;
startscreen[6991] <= 1'b1;
startscreen[6992] <= 1'b1;
startscreen[6997] <= 1'b1;
startscreen[6998] <= 1'b1;
startscreen[7008] <= 1'b1;
startscreen[7009] <= 1'b1;
startscreen[7010] <= 1'b1;
startscreen[7011] <= 1'b1;
startscreen[7012] <= 1'b1;
startscreen[7013] <= 1'b1;
startscreen[7014] <= 1'b1;
startscreen[7015] <= 1'b1;
startscreen[7016] <= 1'b1;
startscreen[7017] <= 1'b1;
startscreen[7018] <= 1'b1;
startscreen[7019] <= 1'b1;
startscreen[7044] <= 1'b1;
startscreen[7045] <= 1'b1;
startscreen[7046] <= 1'b1;
startscreen[7047] <= 1'b1;
startscreen[7066] <= 1'b1;
startscreen[7068] <= 1'b1;
startscreen[7070] <= 1'b1;
startscreen[7071] <= 1'b1;
startscreen[7073] <= 1'b1;
startscreen[7075] <= 1'b1;
startscreen[7087] <= 1'b1;
startscreen[7088] <= 1'b1;
startscreen[7089] <= 1'b1;
startscreen[7090] <= 1'b1;
startscreen[7091] <= 1'b1;
startscreen[7092] <= 1'b1;
startscreen[7094] <= 1'b1;
startscreen[7095] <= 1'b1;
startscreen[7096] <= 1'b1;
startscreen[7097] <= 1'b1;
startscreen[7098] <= 1'b1;
startscreen[7099] <= 1'b1;
startscreen[7110] <= 1'b1;
startscreen[7111] <= 1'b1;
startscreen[7112] <= 1'b1;
startscreen[7113] <= 1'b1;
startscreen[7116] <= 1'b1;
startscreen[7117] <= 1'b1;
startscreen[7118] <= 1'b1;
startscreen[7119] <= 1'b1;
startscreen[7121] <= 1'b1;
startscreen[7123] <= 1'b1;
startscreen[7125] <= 1'b1;
startscreen[7127] <= 1'b1;
startscreen[7128] <= 1'b1;
startscreen[7130] <= 1'b1;
startscreen[7133] <= 1'b1;
startscreen[7134] <= 1'b1;
startscreen[7136] <= 1'b1;
startscreen[7137] <= 1'b1;
startscreen[7147] <= 1'b1;
startscreen[7148] <= 1'b1;
startscreen[7149] <= 1'b1;
startscreen[7150] <= 1'b1;
startscreen[7164] <= 1'b1;
startscreen[7166] <= 1'b1;
startscreen[7173] <= 1'b1;
startscreen[7174] <= 1'b1;
startscreen[7175] <= 1'b1;
startscreen[7176] <= 1'b1;
startscreen[7179] <= 1'b1;
startscreen[7180] <= 1'b1;
startscreen[7181] <= 1'b1;
startscreen[7183] <= 1'b1;
startscreen[7184] <= 1'b1;
startscreen[7185] <= 1'b1;
startscreen[7192] <= 1'b1;
startscreen[7193] <= 1'b1;
startscreen[7195] <= 1'b1;
startscreen[7196] <= 1'b1;
startscreen[7198] <= 1'b1;
startscreen[7199] <= 1'b1;
startscreen[7200] <= 1'b1;
startscreen[7201] <= 1'b1;
startscreen[7203] <= 1'b1;
startscreen[7204] <= 1'b1;
startscreen[7205] <= 1'b1;
startscreen[7215] <= 1'b1;
startscreen[7216] <= 1'b1;
startscreen[7217] <= 1'b1;
startscreen[7218] <= 1'b1;
startscreen[7219] <= 1'b1;
startscreen[7222] <= 1'b1;
startscreen[7223] <= 1'b1;
startscreen[7224] <= 1'b1;
startscreen[7225] <= 1'b1;
startscreen[7227] <= 1'b1;
startscreen[7236] <= 1'b1;
startscreen[7237] <= 1'b1;
startscreen[7238] <= 1'b1;
startscreen[7239] <= 1'b1;
startscreen[7241] <= 1'b1;
startscreen[7242] <= 1'b1;
startscreen[7245] <= 1'b1;
startscreen[7246] <= 1'b1;
startscreen[7247] <= 1'b1;
startscreen[7248] <= 1'b1;
startscreen[7268] <= 1'b1;
startscreen[7269] <= 1'b1;
startscreen[7270] <= 1'b1;
startscreen[7271] <= 1'b1;
startscreen[7272] <= 1'b1;
startscreen[7294] <= 1'b1;
startscreen[7295] <= 1'b1;
startscreen[7296] <= 1'b1;
startscreen[7297] <= 1'b1;
startscreen[7300] <= 1'b1;
startscreen[7303] <= 1'b1;
startscreen[7304] <= 1'b1;
startscreen[7305] <= 1'b1;
startscreen[7307] <= 1'b1;
startscreen[7308] <= 1'b1;
startscreen[7310] <= 1'b1;
startscreen[7311] <= 1'b1;
startscreen[7312] <= 1'b1;
startscreen[7323] <= 1'b1;
startscreen[7324] <= 1'b1;
startscreen[7325] <= 1'b1;
startscreen[7326] <= 1'b1;
startscreen[7327] <= 1'b1;
startscreen[7328] <= 1'b1;
startscreen[7329] <= 1'b1;
startscreen[7331] <= 1'b1;
startscreen[7333] <= 1'b1;
startscreen[7334] <= 1'b1;
startscreen[7335] <= 1'b1;
startscreen[7336] <= 1'b1;
startscreen[7337] <= 1'b1;
startscreen[7350] <= 1'b1;
startscreen[7351] <= 1'b1;
startscreen[7352] <= 1'b1;
startscreen[7353] <= 1'b1;
startscreen[7354] <= 1'b1;
startscreen[7355] <= 1'b1;
startscreen[7356] <= 1'b1;
startscreen[7357] <= 1'b1;
startscreen[7359] <= 1'b1;
startscreen[7360] <= 1'b1;
startscreen[7362] <= 1'b1;
startscreen[7363] <= 1'b1;
startscreen[7372] <= 1'b1;
startscreen[7374] <= 1'b1;
startscreen[7375] <= 1'b1;
startscreen[7376] <= 1'b1;
startscreen[7377] <= 1'b1;
startscreen[7378] <= 1'b1;
startscreen[7379] <= 1'b1;
startscreen[7380] <= 1'b1;
startscreen[7381] <= 1'b1;
startscreen[7383] <= 1'b1;
startscreen[7384] <= 1'b1;
startscreen[7385] <= 1'b1;
startscreen[7404] <= 1'b1;
startscreen[7405] <= 1'b1;
startscreen[7406] <= 1'b1;
startscreen[7409] <= 1'b1;
startscreen[7410] <= 1'b1;
startscreen[7412] <= 1'b1;
startscreen[7413] <= 1'b1;
startscreen[7415] <= 1'b1;
startscreen[7416] <= 1'b1;
startscreen[7418] <= 1'b1;
startscreen[7426] <= 1'b1;
startscreen[7427] <= 1'b1;
startscreen[7428] <= 1'b1;
startscreen[7429] <= 1'b1;
startscreen[7430] <= 1'b1;
startscreen[7431] <= 1'b1;
startscreen[7432] <= 1'b1;
startscreen[7434] <= 1'b1;
startscreen[7436] <= 1'b1;
startscreen[7437] <= 1'b1;
startscreen[7438] <= 1'b1;
startscreen[7439] <= 1'b1;
startscreen[7440] <= 1'b1;
startscreen[7464] <= 1'b1;
startscreen[7465] <= 1'b1;
startscreen[7466] <= 1'b1;
startscreen[7467] <= 1'b1;
startscreen[7468] <= 1'b1;
startscreen[7469] <= 1'b1;
startscreen[7486] <= 1'b1;
startscreen[7487] <= 1'b1;
startscreen[7489] <= 1'b1;
startscreen[7490] <= 1'b1;
startscreen[7491] <= 1'b1;
startscreen[7493] <= 1'b1;
startscreen[7494] <= 1'b1;
startscreen[7497] <= 1'b1;
startscreen[7498] <= 1'b1;
startscreen[7505] <= 1'b1;
startscreen[7506] <= 1'b1;
startscreen[7507] <= 1'b1;
startscreen[7510] <= 1'b1;
startscreen[7511] <= 1'b1;
startscreen[7512] <= 1'b1;
startscreen[7513] <= 1'b1;
startscreen[7514] <= 1'b1;
startscreen[7515] <= 1'b1;
startscreen[7517] <= 1'b1;
startscreen[7518] <= 1'b1;
startscreen[7519] <= 1'b1;
startscreen[7520] <= 1'b1;
startscreen[7530] <= 1'b1;
startscreen[7531] <= 1'b1;
startscreen[7533] <= 1'b1;
startscreen[7535] <= 1'b1;
startscreen[7536] <= 1'b1;
startscreen[7537] <= 1'b1;
startscreen[7538] <= 1'b1;
startscreen[7540] <= 1'b1;
startscreen[7541] <= 1'b1;
startscreen[7543] <= 1'b1;
startscreen[7544] <= 1'b1;
startscreen[7546] <= 1'b1;
startscreen[7547] <= 1'b1;
startscreen[7549] <= 1'b1;
startscreen[7550] <= 1'b1;
startscreen[7552] <= 1'b1;
startscreen[7554] <= 1'b1;
startscreen[7555] <= 1'b1;
startscreen[7557] <= 1'b1;
startscreen[7567] <= 1'b1;
startscreen[7568] <= 1'b1;
startscreen[7569] <= 1'b1;
startscreen[7570] <= 1'b1;
startscreen[7584] <= 1'b1;
startscreen[7586] <= 1'b1;
startscreen[7593] <= 1'b1;
startscreen[7594] <= 1'b1;
startscreen[7595] <= 1'b1;
startscreen[7596] <= 1'b1;
startscreen[7598] <= 1'b1;
startscreen[7599] <= 1'b1;
startscreen[7602] <= 1'b1;
startscreen[7603] <= 1'b1;
startscreen[7604] <= 1'b1;
startscreen[7605] <= 1'b1;
startscreen[7611] <= 1'b1;
startscreen[7614] <= 1'b1;
startscreen[7616] <= 1'b1;
startscreen[7621] <= 1'b1;
startscreen[7622] <= 1'b1;
startscreen[7623] <= 1'b1;
startscreen[7624] <= 1'b1;
startscreen[7625] <= 1'b1;
startscreen[7626] <= 1'b1;
startscreen[7634] <= 1'b1;
startscreen[7635] <= 1'b1;
startscreen[7639] <= 1'b1;
startscreen[7645] <= 1'b1;
startscreen[7646] <= 1'b1;
startscreen[7647] <= 1'b1;
startscreen[7655] <= 1'b1;
startscreen[7656] <= 1'b1;
startscreen[7659] <= 1'b1;
startscreen[7660] <= 1'b1;
startscreen[7666] <= 1'b1;
startscreen[7667] <= 1'b1;
startscreen[7668] <= 1'b1;
startscreen[7689] <= 1'b1;
startscreen[7690] <= 1'b1;
startscreen[7691] <= 1'b1;
startscreen[7692] <= 1'b1;
startscreen[7693] <= 1'b1;
startscreen[7714] <= 1'b1;
startscreen[7715] <= 1'b1;
startscreen[7716] <= 1'b1;
startscreen[7717] <= 1'b1;
startscreen[7719] <= 1'b1;
startscreen[7720] <= 1'b1;
startscreen[7722] <= 1'b1;
startscreen[7723] <= 1'b1;
startscreen[7728] <= 1'b1;
startscreen[7729] <= 1'b1;
startscreen[7733] <= 1'b1;
startscreen[7743] <= 1'b1;
startscreen[7745] <= 1'b1;
startscreen[7746] <= 1'b1;
startscreen[7747] <= 1'b1;
startscreen[7748] <= 1'b1;
startscreen[7753] <= 1'b1;
startscreen[7754] <= 1'b1;
startscreen[7755] <= 1'b1;
startscreen[7756] <= 1'b1;
startscreen[7757] <= 1'b1;
startscreen[7758] <= 1'b1;
startscreen[7769] <= 1'b1;
startscreen[7770] <= 1'b1;
startscreen[7772] <= 1'b1;
startscreen[7773] <= 1'b1;
startscreen[7774] <= 1'b1;
startscreen[7775] <= 1'b1;
startscreen[7780] <= 1'b1;
startscreen[7781] <= 1'b1;
startscreen[7782] <= 1'b1;
startscreen[7783] <= 1'b1;
startscreen[7790] <= 1'b1;
startscreen[7791] <= 1'b1;
startscreen[7792] <= 1'b1;
startscreen[7793] <= 1'b1;
startscreen[7794] <= 1'b1;
startscreen[7795] <= 1'b1;
startscreen[7801] <= 1'b1;
startscreen[7802] <= 1'b1;
startscreen[7803] <= 1'b1;
startscreen[7805] <= 1'b1;
startscreen[7831] <= 1'b1;
startscreen[7832] <= 1'b1;
startscreen[7845] <= 1'b1;
startscreen[7846] <= 1'b1;
startscreen[7847] <= 1'b1;
startscreen[7848] <= 1'b1;
startscreen[7849] <= 1'b1;
startscreen[7850] <= 1'b1;
startscreen[7851] <= 1'b1;
startscreen[7856] <= 1'b1;
startscreen[7857] <= 1'b1;
startscreen[7858] <= 1'b1;
startscreen[7859] <= 1'b1;
startscreen[7860] <= 1'b1;
startscreen[7861] <= 1'b1;
startscreen[7862] <= 1'b1;
startscreen[7885] <= 1'b1;
startscreen[7886] <= 1'b1;
startscreen[7888] <= 1'b1;
startscreen[7889] <= 1'b1;
startscreen[7890] <= 1'b1;
startscreen[7910] <= 1'b1;
startscreen[7911] <= 1'b1;
startscreen[7912] <= 1'b1;
startscreen[7913] <= 1'b1;
startscreen[7925] <= 1'b1;
startscreen[7926] <= 1'b1;
startscreen[7927] <= 1'b1;
startscreen[7928] <= 1'b1;
startscreen[7929] <= 1'b1;
startscreen[7930] <= 1'b1;
startscreen[7931] <= 1'b1;
startscreen[7935] <= 1'b1;
startscreen[7936] <= 1'b1;
startscreen[7937] <= 1'b1;
startscreen[7938] <= 1'b1;
startscreen[7939] <= 1'b1;
startscreen[7940] <= 1'b1;
startscreen[7950] <= 1'b1;
startscreen[7951] <= 1'b1;
startscreen[7952] <= 1'b1;
startscreen[7953] <= 1'b1;
startscreen[7954] <= 1'b1;
startscreen[7955] <= 1'b1;
startscreen[7956] <= 1'b1;
startscreen[7958] <= 1'b1;
startscreen[7960] <= 1'b1;
startscreen[7961] <= 1'b1;
startscreen[7967] <= 1'b1;
startscreen[7968] <= 1'b1;
startscreen[7987] <= 1'b1;
startscreen[7988] <= 1'b1;
startscreen[7989] <= 1'b1;
startscreen[7990] <= 1'b1;
startscreen[8005] <= 1'b1;
startscreen[8006] <= 1'b1;
startscreen[8013] <= 1'b1;
startscreen[8014] <= 1'b1;
startscreen[8015] <= 1'b1;
startscreen[8016] <= 1'b1;
startscreen[8018] <= 1'b1;
startscreen[8019] <= 1'b1;
startscreen[8020] <= 1'b1;
startscreen[8024] <= 1'b1;
startscreen[8025] <= 1'b1;
startscreen[8030] <= 1'b1;
startscreen[8031] <= 1'b1;
startscreen[8033] <= 1'b1;
startscreen[8034] <= 1'b1;
startscreen[8043] <= 1'b1;
startscreen[8045] <= 1'b1;
startscreen[8046] <= 1'b1;
startscreen[8047] <= 1'b1;
startscreen[8054] <= 1'b1;
startscreen[8055] <= 1'b1;
startscreen[8056] <= 1'b1;
startscreen[8057] <= 1'b1;
startscreen[8058] <= 1'b1;
startscreen[8067] <= 1'b1;
startscreen[8075] <= 1'b1;
startscreen[8076] <= 1'b1;
startscreen[8077] <= 1'b1;
startscreen[8078] <= 1'b1;
startscreen[8088] <= 1'b1;
startscreen[8111] <= 1'b1;
startscreen[8112] <= 1'b1;
startscreen[8113] <= 1'b1;
startscreen[8114] <= 1'b1;
startscreen[8134] <= 1'b1;
startscreen[8135] <= 1'b1;
startscreen[8137] <= 1'b1;
startscreen[8139] <= 1'b1;
startscreen[8140] <= 1'b1;
startscreen[8141] <= 1'b1;
startscreen[8150] <= 1'b1;
startscreen[8153] <= 1'b1;
startscreen[8154] <= 1'b1;
startscreen[8163] <= 1'b1;
startscreen[8164] <= 1'b1;
startscreen[8165] <= 1'b1;
startscreen[8175] <= 1'b1;
startscreen[8176] <= 1'b1;
startscreen[8177] <= 1'b1;
startscreen[8178] <= 1'b1;
startscreen[8188] <= 1'b1;
startscreen[8189] <= 1'b1;
startscreen[8190] <= 1'b1;
startscreen[8191] <= 1'b1;
startscreen[8192] <= 1'b1;
startscreen[8202] <= 1'b1;
startscreen[8203] <= 1'b1;
startscreen[8209] <= 1'b1;
startscreen[8210] <= 1'b1;
startscreen[8212] <= 1'b1;
startscreen[8213] <= 1'b1;
startscreen[8214] <= 1'b1;
startscreen[8223] <= 1'b1;
startscreen[8224] <= 1'b1;
startscreen[8225] <= 1'b1;
startscreen[8226] <= 1'b1;
startscreen[8249] <= 1'b1;
startscreen[8250] <= 1'b1;
startscreen[8252] <= 1'b1;
startscreen[8264] <= 1'b1;
startscreen[8265] <= 1'b1;
startscreen[8266] <= 1'b1;
startscreen[8267] <= 1'b1;
startscreen[8268] <= 1'b1;
startscreen[8279] <= 1'b1;
startscreen[8280] <= 1'b1;
startscreen[8281] <= 1'b1;
startscreen[8282] <= 1'b1;
startscreen[8283] <= 1'b1;
startscreen[8306] <= 1'b1;
startscreen[8307] <= 1'b1;
startscreen[8309] <= 1'b1;
startscreen[8310] <= 1'b1;
startscreen[8311] <= 1'b1;
startscreen[8330] <= 1'b1;
startscreen[8332] <= 1'b1;
startscreen[8333] <= 1'b1;
startscreen[8345] <= 1'b1;
startscreen[8346] <= 1'b1;
startscreen[8347] <= 1'b1;
startscreen[8357] <= 1'b1;
startscreen[8358] <= 1'b1;
startscreen[8359] <= 1'b1;
startscreen[8360] <= 1'b1;
startscreen[8361] <= 1'b1;
startscreen[8370] <= 1'b1;
startscreen[8371] <= 1'b1;
startscreen[8372] <= 1'b1;
startscreen[8373] <= 1'b1;
startscreen[8374] <= 1'b1;
startscreen[8375] <= 1'b1;
startscreen[8376] <= 1'b1;
startscreen[8381] <= 1'b1;
startscreen[8387] <= 1'b1;
startscreen[8389] <= 1'b1;
startscreen[8390] <= 1'b1;
startscreen[8407] <= 1'b1;
startscreen[8408] <= 1'b1;
startscreen[8409] <= 1'b1;
startscreen[8410] <= 1'b1;
startscreen[8423] <= 1'b1;
startscreen[8424] <= 1'b1;
startscreen[8425] <= 1'b1;
startscreen[8426] <= 1'b1;
startscreen[8433] <= 1'b1;
startscreen[8434] <= 1'b1;
startscreen[8435] <= 1'b1;
startscreen[8436] <= 1'b1;
startscreen[8437] <= 1'b1;
startscreen[8438] <= 1'b1;
startscreen[8439] <= 1'b1;
startscreen[8450] <= 1'b1;
startscreen[8452] <= 1'b1;
startscreen[8453] <= 1'b1;
startscreen[8464] <= 1'b1;
startscreen[8466] <= 1'b1;
startscreen[8467] <= 1'b1;
startscreen[8473] <= 1'b1;
startscreen[8474] <= 1'b1;
startscreen[8475] <= 1'b1;
startscreen[8476] <= 1'b1;
startscreen[8477] <= 1'b1;
startscreen[8494] <= 1'b1;
startscreen[8495] <= 1'b1;
startscreen[8497] <= 1'b1;
startscreen[8531] <= 1'b1;
startscreen[8532] <= 1'b1;
startscreen[8533] <= 1'b1;
startscreen[8534] <= 1'b1;
startscreen[8536] <= 1'b1;
startscreen[8554] <= 1'b1;
startscreen[8555] <= 1'b1;
startscreen[8556] <= 1'b1;
startscreen[8557] <= 1'b1;
startscreen[8558] <= 1'b1;
startscreen[8559] <= 1'b1;
startscreen[8560] <= 1'b1;
startscreen[8571] <= 1'b1;
startscreen[8572] <= 1'b1;
startscreen[8574] <= 1'b1;
startscreen[8583] <= 1'b1;
startscreen[8595] <= 1'b1;
startscreen[8596] <= 1'b1;
startscreen[8597] <= 1'b1;
startscreen[8598] <= 1'b1;
startscreen[8599] <= 1'b1;
startscreen[8607] <= 1'b1;
startscreen[8608] <= 1'b1;
startscreen[8609] <= 1'b1;
startscreen[8610] <= 1'b1;
startscreen[8611] <= 1'b1;
startscreen[8629] <= 1'b1;
startscreen[8631] <= 1'b1;
startscreen[8632] <= 1'b1;
startscreen[8633] <= 1'b1;
startscreen[8644] <= 1'b1;
startscreen[8645] <= 1'b1;
startscreen[8646] <= 1'b1;
startscreen[8647] <= 1'b1;
startscreen[8669] <= 1'b1;
startscreen[8671] <= 1'b1;
startscreen[8672] <= 1'b1;
startscreen[8683] <= 1'b1;
startscreen[8684] <= 1'b1;
startscreen[8685] <= 1'b1;
startscreen[8686] <= 1'b1;
startscreen[8687] <= 1'b1;
startscreen[8700] <= 1'b1;
startscreen[8701] <= 1'b1;
startscreen[8702] <= 1'b1;
startscreen[8703] <= 1'b1;
startscreen[8727] <= 1'b1;
startscreen[8728] <= 1'b1;
startscreen[8729] <= 1'b1;
startscreen[8731] <= 1'b1;
startscreen[8732] <= 1'b1;
startscreen[8733] <= 1'b1;
startscreen[8750] <= 1'b1;
startscreen[8753] <= 1'b1;
startscreen[8765] <= 1'b1;
startscreen[8766] <= 1'b1;
startscreen[8778] <= 1'b1;
startscreen[8781] <= 1'b1;
startscreen[8790] <= 1'b1;
startscreen[8793] <= 1'b1;
startscreen[8794] <= 1'b1;
startscreen[8795] <= 1'b1;
startscreen[8807] <= 1'b1;
startscreen[8808] <= 1'b1;
startscreen[8810] <= 1'b1;
startscreen[8827] <= 1'b1;
startscreen[8828] <= 1'b1;
startscreen[8829] <= 1'b1;
startscreen[8830] <= 1'b1;
startscreen[8842] <= 1'b1;
startscreen[8844] <= 1'b1;
startscreen[8845] <= 1'b1;
startscreen[8846] <= 1'b1;
startscreen[8853] <= 1'b1;
startscreen[8854] <= 1'b1;
startscreen[8855] <= 1'b1;
startscreen[8856] <= 1'b1;
startscreen[8858] <= 1'b1;
startscreen[8869] <= 1'b1;
startscreen[8870] <= 1'b1;
startscreen[8871] <= 1'b1;
startscreen[8872] <= 1'b1;
startscreen[8873] <= 1'b1;
startscreen[8884] <= 1'b1;
startscreen[8886] <= 1'b1;
startscreen[8887] <= 1'b1;
startscreen[8893] <= 1'b1;
startscreen[8894] <= 1'b1;
startscreen[8895] <= 1'b1;
startscreen[8914] <= 1'b1;
startscreen[8952] <= 1'b1;
startscreen[8953] <= 1'b1;
startscreen[8954] <= 1'b1;
startscreen[8956] <= 1'b1;
startscreen[8958] <= 1'b1;
startscreen[8974] <= 1'b1;
startscreen[8975] <= 1'b1;
startscreen[8976] <= 1'b1;
startscreen[8977] <= 1'b1;
startscreen[8979] <= 1'b1;
startscreen[8992] <= 1'b1;
startscreen[8993] <= 1'b1;
startscreen[8994] <= 1'b1;
startscreen[9016] <= 1'b1;
startscreen[9017] <= 1'b1;
startscreen[9018] <= 1'b1;
startscreen[9019] <= 1'b1;
startscreen[9026] <= 1'b1;
startscreen[9027] <= 1'b1;
startscreen[9029] <= 1'b1;
startscreen[9030] <= 1'b1;
startscreen[9048] <= 1'b1;
startscreen[9049] <= 1'b1;
startscreen[9051] <= 1'b1;
startscreen[9052] <= 1'b1;
startscreen[9064] <= 1'b1;
startscreen[9065] <= 1'b1;
startscreen[9066] <= 1'b1;
startscreen[9067] <= 1'b1;
startscreen[9092] <= 1'b1;
startscreen[9103] <= 1'b1;
startscreen[9104] <= 1'b1;
startscreen[9105] <= 1'b1;
startscreen[9106] <= 1'b1;
startscreen[9121] <= 1'b1;
startscreen[9122] <= 1'b1;
startscreen[9123] <= 1'b1;
startscreen[9124] <= 1'b1;
startscreen[9148] <= 1'b1;
startscreen[9149] <= 1'b1;
startscreen[9150] <= 1'b1;
startscreen[9152] <= 1'b1;
startscreen[9153] <= 1'b1;
startscreen[9154] <= 1'b1;
startscreen[9155] <= 1'b1;
startscreen[9170] <= 1'b1;
startscreen[9171] <= 1'b1;
startscreen[9172] <= 1'b1;
startscreen[9173] <= 1'b1;
startscreen[9198] <= 1'b1;
startscreen[9199] <= 1'b1;
startscreen[9200] <= 1'b1;
startscreen[9201] <= 1'b1;
startscreen[9202] <= 1'b1;
startscreen[9210] <= 1'b1;
startscreen[9212] <= 1'b1;
startscreen[9213] <= 1'b1;
startscreen[9214] <= 1'b1;
startscreen[9227] <= 1'b1;
startscreen[9247] <= 1'b1;
startscreen[9248] <= 1'b1;
startscreen[9249] <= 1'b1;
startscreen[9250] <= 1'b1;
startscreen[9261] <= 1'b1;
startscreen[9263] <= 1'b1;
startscreen[9264] <= 1'b1;
startscreen[9265] <= 1'b1;
startscreen[9273] <= 1'b1;
startscreen[9274] <= 1'b1;
startscreen[9275] <= 1'b1;
startscreen[9276] <= 1'b1;
startscreen[9277] <= 1'b1;
startscreen[9289] <= 1'b1;
startscreen[9290] <= 1'b1;
startscreen[9291] <= 1'b1;
startscreen[9292] <= 1'b1;
startscreen[9305] <= 1'b1;
startscreen[9306] <= 1'b1;
startscreen[9308] <= 1'b1;
startscreen[9313] <= 1'b1;
startscreen[9314] <= 1'b1;
startscreen[9315] <= 1'b1;
startscreen[9316] <= 1'b1;
startscreen[9334] <= 1'b1;
startscreen[9335] <= 1'b1;
startscreen[9336] <= 1'b1;
startscreen[9373] <= 1'b1;
startscreen[9374] <= 1'b1;
startscreen[9375] <= 1'b1;
startscreen[9376] <= 1'b1;
startscreen[9377] <= 1'b1;
startscreen[9378] <= 1'b1;
startscreen[9379] <= 1'b1;
startscreen[9380] <= 1'b1;
startscreen[9394] <= 1'b1;
startscreen[9395] <= 1'b1;
startscreen[9396] <= 1'b1;
startscreen[9397] <= 1'b1;
startscreen[9398] <= 1'b1;
startscreen[9412] <= 1'b1;
startscreen[9414] <= 1'b1;
startscreen[9415] <= 1'b1;
startscreen[9436] <= 1'b1;
startscreen[9437] <= 1'b1;
startscreen[9438] <= 1'b1;
startscreen[9439] <= 1'b1;
startscreen[9446] <= 1'b1;
startscreen[9448] <= 1'b1;
startscreen[9449] <= 1'b1;
startscreen[9468] <= 1'b1;
startscreen[9469] <= 1'b1;
startscreen[9470] <= 1'b1;
startscreen[9471] <= 1'b1;
startscreen[9485] <= 1'b1;
startscreen[9486] <= 1'b1;
startscreen[9487] <= 1'b1;
startscreen[9509] <= 1'b1;
startscreen[9511] <= 1'b1;
startscreen[9512] <= 1'b1;
startscreen[9522] <= 1'b1;
startscreen[9523] <= 1'b1;
startscreen[9524] <= 1'b1;
startscreen[9525] <= 1'b1;
startscreen[9526] <= 1'b1;
startscreen[9541] <= 1'b1;
startscreen[9542] <= 1'b1;
startscreen[9543] <= 1'b1;
startscreen[9544] <= 1'b1;
startscreen[9569] <= 1'b1;
startscreen[9570] <= 1'b1;
startscreen[9571] <= 1'b1;
startscreen[9572] <= 1'b1;
startscreen[9573] <= 1'b1;
startscreen[9574] <= 1'b1;
startscreen[9575] <= 1'b1;
startscreen[9576] <= 1'b1;
startscreen[9590] <= 1'b1;
startscreen[9592] <= 1'b1;
startscreen[9593] <= 1'b1;
startscreen[9619] <= 1'b1;
startscreen[9621] <= 1'b1;
startscreen[9622] <= 1'b1;
startscreen[9631] <= 1'b1;
startscreen[9633] <= 1'b1;
startscreen[9647] <= 1'b1;
startscreen[9648] <= 1'b1;
startscreen[9667] <= 1'b1;
startscreen[9668] <= 1'b1;
startscreen[9669] <= 1'b1;
startscreen[9670] <= 1'b1;
startscreen[9679] <= 1'b1;
startscreen[9681] <= 1'b1;
startscreen[9682] <= 1'b1;
startscreen[9684] <= 1'b1;
startscreen[9693] <= 1'b1;
startscreen[9694] <= 1'b1;
startscreen[9695] <= 1'b1;
startscreen[9696] <= 1'b1;
startscreen[9708] <= 1'b1;
startscreen[9709] <= 1'b1;
startscreen[9710] <= 1'b1;
startscreen[9725] <= 1'b1;
startscreen[9726] <= 1'b1;
startscreen[9728] <= 1'b1;
startscreen[9733] <= 1'b1;
startscreen[9734] <= 1'b1;
startscreen[9735] <= 1'b1;
startscreen[9736] <= 1'b1;
startscreen[9737] <= 1'b1;
startscreen[9754] <= 1'b1;
startscreen[9756] <= 1'b1;
startscreen[9757] <= 1'b1;
startscreen[9795] <= 1'b1;
startscreen[9796] <= 1'b1;
startscreen[9798] <= 1'b1;
startscreen[9801] <= 1'b1;
startscreen[9802] <= 1'b1;
startscreen[9814] <= 1'b1;
startscreen[9815] <= 1'b1;
startscreen[9817] <= 1'b1;
startscreen[9832] <= 1'b1;
startscreen[9834] <= 1'b1;
startscreen[9835] <= 1'b1;
startscreen[9856] <= 1'b1;
startscreen[9857] <= 1'b1;
startscreen[9858] <= 1'b1;
startscreen[9859] <= 1'b1;
startscreen[9865] <= 1'b1;
startscreen[9866] <= 1'b1;
startscreen[9868] <= 1'b1;
startscreen[9887] <= 1'b1;
startscreen[9888] <= 1'b1;
startscreen[9889] <= 1'b1;
startscreen[9890] <= 1'b1;
startscreen[9905] <= 1'b1;
startscreen[9906] <= 1'b1;
startscreen[9907] <= 1'b1;
startscreen[9908] <= 1'b1;
startscreen[9930] <= 1'b1;
startscreen[9931] <= 1'b1;
startscreen[9932] <= 1'b1;
startscreen[9942] <= 1'b1;
startscreen[9943] <= 1'b1;
startscreen[9944] <= 1'b1;
startscreen[9945] <= 1'b1;
startscreen[9946] <= 1'b1;
startscreen[9961] <= 1'b1;
startscreen[9962] <= 1'b1;
startscreen[9964] <= 1'b1;
startscreen[9965] <= 1'b1;
startscreen[9993] <= 1'b1;
startscreen[9995] <= 1'b1;
startscreen[9996] <= 1'b1;
startscreen[9997] <= 1'b1;
startscreen[9998] <= 1'b1;
startscreen[10010] <= 1'b1;
startscreen[10011] <= 1'b1;
startscreen[10012] <= 1'b1;
startscreen[10013] <= 1'b1;
startscreen[10039] <= 1'b1;
startscreen[10040] <= 1'b1;
startscreen[10041] <= 1'b1;
startscreen[10042] <= 1'b1;
startscreen[10052] <= 1'b1;
startscreen[10053] <= 1'b1;
startscreen[10067] <= 1'b1;
startscreen[10068] <= 1'b1;
startscreen[10069] <= 1'b1;
startscreen[10087] <= 1'b1;
startscreen[10088] <= 1'b1;
startscreen[10089] <= 1'b1;
startscreen[10090] <= 1'b1;
startscreen[10091] <= 1'b1;
startscreen[10092] <= 1'b1;
startscreen[10093] <= 1'b1;
startscreen[10096] <= 1'b1;
startscreen[10099] <= 1'b1;
startscreen[10100] <= 1'b1;
startscreen[10103] <= 1'b1;
startscreen[10113] <= 1'b1;
startscreen[10114] <= 1'b1;
startscreen[10115] <= 1'b1;
startscreen[10116] <= 1'b1;
startscreen[10128] <= 1'b1;
startscreen[10129] <= 1'b1;
startscreen[10130] <= 1'b1;
startscreen[10131] <= 1'b1;
startscreen[10145] <= 1'b1;
startscreen[10146] <= 1'b1;
startscreen[10148] <= 1'b1;
startscreen[10154] <= 1'b1;
startscreen[10155] <= 1'b1;
startscreen[10157] <= 1'b1;
startscreen[10158] <= 1'b1;
startscreen[10175] <= 1'b1;
startscreen[10176] <= 1'b1;
startscreen[10178] <= 1'b1;
startscreen[10217] <= 1'b1;
startscreen[10220] <= 1'b1;
startscreen[10234] <= 1'b1;
startscreen[10235] <= 1'b1;
startscreen[10237] <= 1'b1;
startscreen[10253] <= 1'b1;
startscreen[10254] <= 1'b1;
startscreen[10255] <= 1'b1;
startscreen[10256] <= 1'b1;
startscreen[10272] <= 1'b1;
startscreen[10273] <= 1'b1;
startscreen[10274] <= 1'b1;
startscreen[10275] <= 1'b1;
startscreen[10276] <= 1'b1;
startscreen[10277] <= 1'b1;
startscreen[10278] <= 1'b1;
startscreen[10279] <= 1'b1;
startscreen[10285] <= 1'b1;
startscreen[10286] <= 1'b1;
startscreen[10287] <= 1'b1;
startscreen[10288] <= 1'b1;
startscreen[10307] <= 1'b1;
startscreen[10308] <= 1'b1;
startscreen[10309] <= 1'b1;
startscreen[10325] <= 1'b1;
startscreen[10327] <= 1'b1;
startscreen[10328] <= 1'b1;
startscreen[10350] <= 1'b1;
startscreen[10351] <= 1'b1;
startscreen[10352] <= 1'b1;
startscreen[10362] <= 1'b1;
startscreen[10363] <= 1'b1;
startscreen[10364] <= 1'b1;
startscreen[10365] <= 1'b1;
startscreen[10382] <= 1'b1;
startscreen[10383] <= 1'b1;
startscreen[10384] <= 1'b1;
startscreen[10385] <= 1'b1;
startscreen[10413] <= 1'b1;
startscreen[10414] <= 1'b1;
startscreen[10416] <= 1'b1;
startscreen[10417] <= 1'b1;
startscreen[10418] <= 1'b1;
startscreen[10419] <= 1'b1;
startscreen[10420] <= 1'b1;
startscreen[10430] <= 1'b1;
startscreen[10431] <= 1'b1;
startscreen[10432] <= 1'b1;
startscreen[10433] <= 1'b1;
startscreen[10452] <= 1'b1;
startscreen[10453] <= 1'b1;
startscreen[10454] <= 1'b1;
startscreen[10455] <= 1'b1;
startscreen[10456] <= 1'b1;
startscreen[10457] <= 1'b1;
startscreen[10460] <= 1'b1;
startscreen[10461] <= 1'b1;
startscreen[10462] <= 1'b1;
startscreen[10470] <= 1'b1;
startscreen[10471] <= 1'b1;
startscreen[10473] <= 1'b1;
startscreen[10487] <= 1'b1;
startscreen[10488] <= 1'b1;
startscreen[10489] <= 1'b1;
startscreen[10507] <= 1'b1;
startscreen[10508] <= 1'b1;
startscreen[10509] <= 1'b1;
startscreen[10510] <= 1'b1;
startscreen[10511] <= 1'b1;
startscreen[10513] <= 1'b1;
startscreen[10514] <= 1'b1;
startscreen[10515] <= 1'b1;
startscreen[10517] <= 1'b1;
startscreen[10518] <= 1'b1;
startscreen[10520] <= 1'b1;
startscreen[10522] <= 1'b1;
startscreen[10533] <= 1'b1;
startscreen[10534] <= 1'b1;
startscreen[10535] <= 1'b1;
startscreen[10536] <= 1'b1;
startscreen[10548] <= 1'b1;
startscreen[10549] <= 1'b1;
startscreen[10550] <= 1'b1;
startscreen[10551] <= 1'b1;
startscreen[10552] <= 1'b1;
startscreen[10553] <= 1'b1;
startscreen[10554] <= 1'b1;
startscreen[10555] <= 1'b1;
startscreen[10556] <= 1'b1;
startscreen[10557] <= 1'b1;
startscreen[10558] <= 1'b1;
startscreen[10559] <= 1'b1;
startscreen[10560] <= 1'b1;
startscreen[10561] <= 1'b1;
startscreen[10562] <= 1'b1;
startscreen[10563] <= 1'b1;
startscreen[10564] <= 1'b1;
startscreen[10565] <= 1'b1;
startscreen[10566] <= 1'b1;
startscreen[10567] <= 1'b1;
startscreen[10568] <= 1'b1;
startscreen[10569] <= 1'b1;
startscreen[10575] <= 1'b1;
startscreen[10576] <= 1'b1;
startscreen[10577] <= 1'b1;
startscreen[10578] <= 1'b1;
startscreen[10580] <= 1'b1;
startscreen[10581] <= 1'b1;
startscreen[10596] <= 1'b1;
startscreen[10597] <= 1'b1;
startscreen[10598] <= 1'b1;
startscreen[10600] <= 1'b1;
startscreen[10639] <= 1'b1;
startscreen[10640] <= 1'b1;
startscreen[10641] <= 1'b1;
startscreen[10643] <= 1'b1;
startscreen[10654] <= 1'b1;
startscreen[10655] <= 1'b1;
startscreen[10656] <= 1'b1;
startscreen[10657] <= 1'b1;
startscreen[10673] <= 1'b1;
startscreen[10675] <= 1'b1;
startscreen[10676] <= 1'b1;
startscreen[10687] <= 1'b1;
startscreen[10688] <= 1'b1;
startscreen[10689] <= 1'b1;
startscreen[10690] <= 1'b1;
startscreen[10691] <= 1'b1;
startscreen[10692] <= 1'b1;
startscreen[10693] <= 1'b1;
startscreen[10694] <= 1'b1;
startscreen[10696] <= 1'b1;
startscreen[10698] <= 1'b1;
startscreen[10699] <= 1'b1;
startscreen[10705] <= 1'b1;
startscreen[10706] <= 1'b1;
startscreen[10708] <= 1'b1;
startscreen[10727] <= 1'b1;
startscreen[10728] <= 1'b1;
startscreen[10729] <= 1'b1;
startscreen[10730] <= 1'b1;
startscreen[10731] <= 1'b1;
startscreen[10732] <= 1'b1;
startscreen[10734] <= 1'b1;
startscreen[10736] <= 1'b1;
startscreen[10737] <= 1'b1;
startscreen[10738] <= 1'b1;
startscreen[10739] <= 1'b1;
startscreen[10740] <= 1'b1;
startscreen[10741] <= 1'b1;
startscreen[10742] <= 1'b1;
startscreen[10743] <= 1'b1;
startscreen[10745] <= 1'b1;
startscreen[10746] <= 1'b1;
startscreen[10747] <= 1'b1;
startscreen[10748] <= 1'b1;
startscreen[10770] <= 1'b1;
startscreen[10771] <= 1'b1;
startscreen[10772] <= 1'b1;
startscreen[10782] <= 1'b1;
startscreen[10785] <= 1'b1;
startscreen[10802] <= 1'b1;
startscreen[10804] <= 1'b1;
startscreen[10805] <= 1'b1;
startscreen[10834] <= 1'b1;
startscreen[10835] <= 1'b1;
startscreen[10836] <= 1'b1;
startscreen[10837] <= 1'b1;
startscreen[10839] <= 1'b1;
startscreen[10840] <= 1'b1;
startscreen[10841] <= 1'b1;
startscreen[10850] <= 1'b1;
startscreen[10851] <= 1'b1;
startscreen[10852] <= 1'b1;
startscreen[10853] <= 1'b1;
startscreen[10869] <= 1'b1;
startscreen[10870] <= 1'b1;
startscreen[10871] <= 1'b1;
startscreen[10872] <= 1'b1;
startscreen[10874] <= 1'b1;
startscreen[10875] <= 1'b1;
startscreen[10876] <= 1'b1;
startscreen[10877] <= 1'b1;
startscreen[10878] <= 1'b1;
startscreen[10880] <= 1'b1;
startscreen[10881] <= 1'b1;
startscreen[10882] <= 1'b1;
startscreen[10890] <= 1'b1;
startscreen[10891] <= 1'b1;
startscreen[10893] <= 1'b1;
startscreen[10907] <= 1'b1;
startscreen[10908] <= 1'b1;
startscreen[10909] <= 1'b1;
startscreen[10927] <= 1'b1;
startscreen[10928] <= 1'b1;
startscreen[10929] <= 1'b1;
startscreen[10930] <= 1'b1;
startscreen[10932] <= 1'b1;
startscreen[10933] <= 1'b1;
startscreen[10935] <= 1'b1;
startscreen[10940] <= 1'b1;
startscreen[10953] <= 1'b1;
startscreen[10954] <= 1'b1;
startscreen[10955] <= 1'b1;
startscreen[10956] <= 1'b1;
startscreen[10968] <= 1'b1;
startscreen[10969] <= 1'b1;
startscreen[10970] <= 1'b1;
startscreen[10971] <= 1'b1;
startscreen[10973] <= 1'b1;
startscreen[10974] <= 1'b1;
startscreen[10976] <= 1'b1;
startscreen[10977] <= 1'b1;
startscreen[10978] <= 1'b1;
startscreen[10979] <= 1'b1;
startscreen[10980] <= 1'b1;
startscreen[10981] <= 1'b1;
startscreen[10982] <= 1'b1;
startscreen[10988] <= 1'b1;
startscreen[10989] <= 1'b1;
startscreen[10996] <= 1'b1;
startscreen[10998] <= 1'b1;
startscreen[10999] <= 1'b1;
startscreen[11000] <= 1'b1;
startscreen[11001] <= 1'b1;
startscreen[11002] <= 1'b1;
startscreen[11003] <= 1'b1;
startscreen[11017] <= 1'b1;
startscreen[11019] <= 1'b1;
startscreen[11020] <= 1'b1;
startscreen[11023] <= 1'b1;
startscreen[11061] <= 1'b1;
startscreen[11062] <= 1'b1;
startscreen[11064] <= 1'b1;
startscreen[11074] <= 1'b1;
startscreen[11075] <= 1'b1;
startscreen[11076] <= 1'b1;
startscreen[11077] <= 1'b1;
startscreen[11093] <= 1'b1;
startscreen[11095] <= 1'b1;
startscreen[11096] <= 1'b1;
startscreen[11104] <= 1'b1;
startscreen[11105] <= 1'b1;
startscreen[11106] <= 1'b1;
startscreen[11107] <= 1'b1;
startscreen[11108] <= 1'b1;
startscreen[11109] <= 1'b1;
startscreen[11110] <= 1'b1;
startscreen[11111] <= 1'b1;
startscreen[11114] <= 1'b1;
startscreen[11115] <= 1'b1;
startscreen[11116] <= 1'b1;
startscreen[11117] <= 1'b1;
startscreen[11118] <= 1'b1;
startscreen[11119] <= 1'b1;
startscreen[11125] <= 1'b1;
startscreen[11127] <= 1'b1;
startscreen[11128] <= 1'b1;
startscreen[11147] <= 1'b1;
startscreen[11148] <= 1'b1;
startscreen[11149] <= 1'b1;
startscreen[11151] <= 1'b1;
startscreen[11153] <= 1'b1;
startscreen[11155] <= 1'b1;
startscreen[11156] <= 1'b1;
startscreen[11157] <= 1'b1;
startscreen[11158] <= 1'b1;
startscreen[11159] <= 1'b1;
startscreen[11160] <= 1'b1;
startscreen[11161] <= 1'b1;
startscreen[11162] <= 1'b1;
startscreen[11163] <= 1'b1;
startscreen[11165] <= 1'b1;
startscreen[11166] <= 1'b1;
startscreen[11167] <= 1'b1;
startscreen[11168] <= 1'b1;
startscreen[11190] <= 1'b1;
startscreen[11191] <= 1'b1;
startscreen[11192] <= 1'b1;
startscreen[11202] <= 1'b1;
startscreen[11205] <= 1'b1;
startscreen[11222] <= 1'b1;
startscreen[11223] <= 1'b1;
startscreen[11224] <= 1'b1;
startscreen[11225] <= 1'b1;
startscreen[11257] <= 1'b1;
startscreen[11258] <= 1'b1;
startscreen[11259] <= 1'b1;
startscreen[11260] <= 1'b1;
startscreen[11261] <= 1'b1;
startscreen[11262] <= 1'b1;
startscreen[11270] <= 1'b1;
startscreen[11271] <= 1'b1;
startscreen[11272] <= 1'b1;
startscreen[11273] <= 1'b1;
startscreen[11286] <= 1'b1;
startscreen[11287] <= 1'b1;
startscreen[11288] <= 1'b1;
startscreen[11289] <= 1'b1;
startscreen[11290] <= 1'b1;
startscreen[11292] <= 1'b1;
startscreen[11293] <= 1'b1;
startscreen[11294] <= 1'b1;
startscreen[11295] <= 1'b1;
startscreen[11297] <= 1'b1;
startscreen[11298] <= 1'b1;
startscreen[11299] <= 1'b1;
startscreen[11300] <= 1'b1;
startscreen[11301] <= 1'b1;
startscreen[11302] <= 1'b1;
startscreen[11312] <= 1'b1;
startscreen[11313] <= 1'b1;
startscreen[11327] <= 1'b1;
startscreen[11328] <= 1'b1;
startscreen[11329] <= 1'b1;
startscreen[11347] <= 1'b1;
startscreen[11348] <= 1'b1;
startscreen[11349] <= 1'b1;
startscreen[11350] <= 1'b1;
startscreen[11351] <= 1'b1;
startscreen[11352] <= 1'b1;
startscreen[11353] <= 1'b1;
startscreen[11354] <= 1'b1;
startscreen[11355] <= 1'b1;
startscreen[11356] <= 1'b1;
startscreen[11357] <= 1'b1;
startscreen[11373] <= 1'b1;
startscreen[11374] <= 1'b1;
startscreen[11375] <= 1'b1;
startscreen[11376] <= 1'b1;
startscreen[11388] <= 1'b1;
startscreen[11389] <= 1'b1;
startscreen[11390] <= 1'b1;
startscreen[11391] <= 1'b1;
startscreen[11392] <= 1'b1;
startscreen[11393] <= 1'b1;
startscreen[11394] <= 1'b1;
startscreen[11395] <= 1'b1;
startscreen[11397] <= 1'b1;
startscreen[11398] <= 1'b1;
startscreen[11400] <= 1'b1;
startscreen[11402] <= 1'b1;
startscreen[11403] <= 1'b1;
startscreen[11404] <= 1'b1;
startscreen[11405] <= 1'b1;
startscreen[11406] <= 1'b1;
startscreen[11407] <= 1'b1;
startscreen[11408] <= 1'b1;
startscreen[11409] <= 1'b1;
startscreen[11417] <= 1'b1;
startscreen[11421] <= 1'b1;
startscreen[11422] <= 1'b1;
startscreen[11423] <= 1'b1;
startscreen[11424] <= 1'b1;
startscreen[11425] <= 1'b1;
startscreen[11438] <= 1'b1;
startscreen[11441] <= 1'b1;
startscreen[11445] <= 1'b1;
startscreen[11482] <= 1'b1;
startscreen[11483] <= 1'b1;
startscreen[11485] <= 1'b1;
startscreen[11486] <= 1'b1;
startscreen[11494] <= 1'b1;
startscreen[11495] <= 1'b1;
startscreen[11496] <= 1'b1;
startscreen[11497] <= 1'b1;
startscreen[11513] <= 1'b1;
startscreen[11514] <= 1'b1;
startscreen[11515] <= 1'b1;
startscreen[11516] <= 1'b1;
startscreen[11523] <= 1'b1;
startscreen[11524] <= 1'b1;
startscreen[11525] <= 1'b1;
startscreen[11526] <= 1'b1;
startscreen[11527] <= 1'b1;
startscreen[11528] <= 1'b1;
startscreen[11529] <= 1'b1;
startscreen[11530] <= 1'b1;
startscreen[11531] <= 1'b1;
startscreen[11532] <= 1'b1;
startscreen[11536] <= 1'b1;
startscreen[11538] <= 1'b1;
startscreen[11539] <= 1'b1;
startscreen[11545] <= 1'b1;
startscreen[11546] <= 1'b1;
startscreen[11547] <= 1'b1;
startscreen[11548] <= 1'b1;
startscreen[11567] <= 1'b1;
startscreen[11568] <= 1'b1;
startscreen[11569] <= 1'b1;
startscreen[11571] <= 1'b1;
startscreen[11573] <= 1'b1;
startscreen[11574] <= 1'b1;
startscreen[11576] <= 1'b1;
startscreen[11577] <= 1'b1;
startscreen[11578] <= 1'b1;
startscreen[11579] <= 1'b1;
startscreen[11580] <= 1'b1;
startscreen[11581] <= 1'b1;
startscreen[11582] <= 1'b1;
startscreen[11583] <= 1'b1;
startscreen[11584] <= 1'b1;
startscreen[11585] <= 1'b1;
startscreen[11586] <= 1'b1;
startscreen[11587] <= 1'b1;
startscreen[11588] <= 1'b1;
startscreen[11610] <= 1'b1;
startscreen[11611] <= 1'b1;
startscreen[11612] <= 1'b1;
startscreen[11622] <= 1'b1;
startscreen[11623] <= 1'b1;
startscreen[11624] <= 1'b1;
startscreen[11625] <= 1'b1;
startscreen[11642] <= 1'b1;
startscreen[11643] <= 1'b1;
startscreen[11644] <= 1'b1;
startscreen[11645] <= 1'b1;
startscreen[11678] <= 1'b1;
startscreen[11679] <= 1'b1;
startscreen[11681] <= 1'b1;
startscreen[11682] <= 1'b1;
startscreen[11690] <= 1'b1;
startscreen[11691] <= 1'b1;
startscreen[11692] <= 1'b1;
startscreen[11693] <= 1'b1;
startscreen[11705] <= 1'b1;
startscreen[11706] <= 1'b1;
startscreen[11707] <= 1'b1;
startscreen[11709] <= 1'b1;
startscreen[11710] <= 1'b1;
startscreen[11711] <= 1'b1;
startscreen[11712] <= 1'b1;
startscreen[11713] <= 1'b1;
startscreen[11720] <= 1'b1;
startscreen[11721] <= 1'b1;
startscreen[11722] <= 1'b1;
startscreen[11730] <= 1'b1;
startscreen[11732] <= 1'b1;
startscreen[11733] <= 1'b1;
startscreen[11747] <= 1'b1;
startscreen[11748] <= 1'b1;
startscreen[11749] <= 1'b1;
startscreen[11767] <= 1'b1;
startscreen[11768] <= 1'b1;
startscreen[11769] <= 1'b1;
startscreen[11770] <= 1'b1;
startscreen[11793] <= 1'b1;
startscreen[11794] <= 1'b1;
startscreen[11795] <= 1'b1;
startscreen[11796] <= 1'b1;
startscreen[11808] <= 1'b1;
startscreen[11809] <= 1'b1;
startscreen[11810] <= 1'b1;
startscreen[11811] <= 1'b1;
startscreen[11839] <= 1'b1;
startscreen[11840] <= 1'b1;
startscreen[11841] <= 1'b1;
startscreen[11845] <= 1'b1;
startscreen[11846] <= 1'b1;
startscreen[11860] <= 1'b1;
startscreen[11861] <= 1'b1;
startscreen[11863] <= 1'b1;
startscreen[11864] <= 1'b1;
startscreen[11867] <= 1'b1;
startscreen[11903] <= 1'b1;
startscreen[11906] <= 1'b1;
startscreen[11907] <= 1'b1;
startscreen[11914] <= 1'b1;
startscreen[11915] <= 1'b1;
startscreen[11916] <= 1'b1;
startscreen[11917] <= 1'b1;
startscreen[11933] <= 1'b1;
startscreen[11935] <= 1'b1;
startscreen[11936] <= 1'b1;
startscreen[11942] <= 1'b1;
startscreen[11943] <= 1'b1;
startscreen[11944] <= 1'b1;
startscreen[11945] <= 1'b1;
startscreen[11946] <= 1'b1;
startscreen[11947] <= 1'b1;
startscreen[11956] <= 1'b1;
startscreen[11957] <= 1'b1;
startscreen[11959] <= 1'b1;
startscreen[11965] <= 1'b1;
startscreen[11966] <= 1'b1;
startscreen[11968] <= 1'b1;
startscreen[11987] <= 1'b1;
startscreen[11988] <= 1'b1;
startscreen[11990] <= 1'b1;
startscreen[12030] <= 1'b1;
startscreen[12031] <= 1'b1;
startscreen[12032] <= 1'b1;
startscreen[12042] <= 1'b1;
startscreen[12043] <= 1'b1;
startscreen[12045] <= 1'b1;
startscreen[12062] <= 1'b1;
startscreen[12063] <= 1'b1;
startscreen[12064] <= 1'b1;
startscreen[12065] <= 1'b1;
startscreen[12099] <= 1'b1;
startscreen[12100] <= 1'b1;
startscreen[12101] <= 1'b1;
startscreen[12102] <= 1'b1;
startscreen[12103] <= 1'b1;
startscreen[12110] <= 1'b1;
startscreen[12111] <= 1'b1;
startscreen[12112] <= 1'b1;
startscreen[12113] <= 1'b1;
startscreen[12125] <= 1'b1;
startscreen[12126] <= 1'b1;
startscreen[12127] <= 1'b1;
startscreen[12128] <= 1'b1;
startscreen[12129] <= 1'b1;
startscreen[12140] <= 1'b1;
startscreen[12142] <= 1'b1;
startscreen[12150] <= 1'b1;
startscreen[12151] <= 1'b1;
startscreen[12152] <= 1'b1;
startscreen[12153] <= 1'b1;
startscreen[12167] <= 1'b1;
startscreen[12168] <= 1'b1;
startscreen[12169] <= 1'b1;
startscreen[12187] <= 1'b1;
startscreen[12188] <= 1'b1;
startscreen[12189] <= 1'b1;
startscreen[12190] <= 1'b1;
startscreen[12213] <= 1'b1;
startscreen[12214] <= 1'b1;
startscreen[12215] <= 1'b1;
startscreen[12216] <= 1'b1;
startscreen[12228] <= 1'b1;
startscreen[12229] <= 1'b1;
startscreen[12230] <= 1'b1;
startscreen[12231] <= 1'b1;
startscreen[12262] <= 1'b1;
startscreen[12263] <= 1'b1;
startscreen[12264] <= 1'b1;
startscreen[12265] <= 1'b1;
startscreen[12266] <= 1'b1;
startscreen[12267] <= 1'b1;
startscreen[12282] <= 1'b1;
startscreen[12283] <= 1'b1;
startscreen[12284] <= 1'b1;
startscreen[12285] <= 1'b1;
startscreen[12286] <= 1'b1;
startscreen[12287] <= 1'b1;
startscreen[12288] <= 1'b1;
startscreen[12324] <= 1'b1;
startscreen[12325] <= 1'b1;
startscreen[12327] <= 1'b1;
startscreen[12334] <= 1'b1;
startscreen[12335] <= 1'b1;
startscreen[12337] <= 1'b1;
startscreen[12353] <= 1'b1;
startscreen[12355] <= 1'b1;
startscreen[12356] <= 1'b1;
startscreen[12361] <= 1'b1;
startscreen[12362] <= 1'b1;
startscreen[12364] <= 1'b1;
startscreen[12365] <= 1'b1;
startscreen[12376] <= 1'b1;
startscreen[12377] <= 1'b1;
startscreen[12378] <= 1'b1;
startscreen[12379] <= 1'b1;
startscreen[12385] <= 1'b1;
startscreen[12386] <= 1'b1;
startscreen[12387] <= 1'b1;
startscreen[12388] <= 1'b1;
startscreen[12407] <= 1'b1;
startscreen[12408] <= 1'b1;
startscreen[12409] <= 1'b1;
startscreen[12450] <= 1'b1;
startscreen[12451] <= 1'b1;
startscreen[12452] <= 1'b1;
startscreen[12462] <= 1'b1;
startscreen[12463] <= 1'b1;
startscreen[12465] <= 1'b1;
startscreen[12482] <= 1'b1;
startscreen[12483] <= 1'b1;
startscreen[12484] <= 1'b1;
startscreen[12485] <= 1'b1;
startscreen[12520] <= 1'b1;
startscreen[12521] <= 1'b1;
startscreen[12522] <= 1'b1;
startscreen[12523] <= 1'b1;
startscreen[12530] <= 1'b1;
startscreen[12531] <= 1'b1;
startscreen[12532] <= 1'b1;
startscreen[12533] <= 1'b1;
startscreen[12544] <= 1'b1;
startscreen[12545] <= 1'b1;
startscreen[12547] <= 1'b1;
startscreen[12548] <= 1'b1;
startscreen[12559] <= 1'b1;
startscreen[12560] <= 1'b1;
startscreen[12561] <= 1'b1;
startscreen[12562] <= 1'b1;
startscreen[12571] <= 1'b1;
startscreen[12572] <= 1'b1;
startscreen[12573] <= 1'b1;
startscreen[12587] <= 1'b1;
startscreen[12588] <= 1'b1;
startscreen[12589] <= 1'b1;
startscreen[12607] <= 1'b1;
startscreen[12608] <= 1'b1;
startscreen[12609] <= 1'b1;
startscreen[12610] <= 1'b1;
startscreen[12633] <= 1'b1;
startscreen[12634] <= 1'b1;
startscreen[12635] <= 1'b1;
startscreen[12636] <= 1'b1;
startscreen[12648] <= 1'b1;
startscreen[12649] <= 1'b1;
startscreen[12650] <= 1'b1;
startscreen[12651] <= 1'b1;
startscreen[12683] <= 1'b1;
startscreen[12684] <= 1'b1;
startscreen[12685] <= 1'b1;
startscreen[12686] <= 1'b1;
startscreen[12687] <= 1'b1;
startscreen[12688] <= 1'b1;
startscreen[12704] <= 1'b1;
startscreen[12705] <= 1'b1;
startscreen[12706] <= 1'b1;
startscreen[12707] <= 1'b1;
startscreen[12744] <= 1'b1;
startscreen[12746] <= 1'b1;
startscreen[12747] <= 1'b1;
startscreen[12754] <= 1'b1;
startscreen[12755] <= 1'b1;
startscreen[12756] <= 1'b1;
startscreen[12757] <= 1'b1;
startscreen[12772] <= 1'b1;
startscreen[12774] <= 1'b1;
startscreen[12775] <= 1'b1;
startscreen[12776] <= 1'b1;
startscreen[12781] <= 1'b1;
startscreen[12782] <= 1'b1;
startscreen[12784] <= 1'b1;
startscreen[12796] <= 1'b1;
startscreen[12798] <= 1'b1;
startscreen[12799] <= 1'b1;
startscreen[12805] <= 1'b1;
startscreen[12807] <= 1'b1;
startscreen[12808] <= 1'b1;
startscreen[12827] <= 1'b1;
startscreen[12828] <= 1'b1;
startscreen[12830] <= 1'b1;
startscreen[12870] <= 1'b1;
startscreen[12871] <= 1'b1;
startscreen[12872] <= 1'b1;
startscreen[12882] <= 1'b1;
startscreen[12884] <= 1'b1;
startscreen[12885] <= 1'b1;
startscreen[12902] <= 1'b1;
startscreen[12904] <= 1'b1;
startscreen[12905] <= 1'b1;
startscreen[12940] <= 1'b1;
startscreen[12941] <= 1'b1;
startscreen[12942] <= 1'b1;
startscreen[12943] <= 1'b1;
startscreen[12950] <= 1'b1;
startscreen[12951] <= 1'b1;
startscreen[12952] <= 1'b1;
startscreen[12953] <= 1'b1;
startscreen[12963] <= 1'b1;
startscreen[12964] <= 1'b1;
startscreen[12965] <= 1'b1;
startscreen[12966] <= 1'b1;
startscreen[12967] <= 1'b1;
startscreen[12979] <= 1'b1;
startscreen[12980] <= 1'b1;
startscreen[12981] <= 1'b1;
startscreen[12982] <= 1'b1;
startscreen[12990] <= 1'b1;
startscreen[12993] <= 1'b1;
startscreen[13007] <= 1'b1;
startscreen[13008] <= 1'b1;
startscreen[13009] <= 1'b1;
startscreen[13027] <= 1'b1;
startscreen[13028] <= 1'b1;
startscreen[13029] <= 1'b1;
startscreen[13030] <= 1'b1;
startscreen[13053] <= 1'b1;
startscreen[13054] <= 1'b1;
startscreen[13055] <= 1'b1;
startscreen[13056] <= 1'b1;
startscreen[13068] <= 1'b1;
startscreen[13069] <= 1'b1;
startscreen[13071] <= 1'b1;
startscreen[13072] <= 1'b1;
startscreen[13105] <= 1'b1;
startscreen[13106] <= 1'b1;
startscreen[13107] <= 1'b1;
startscreen[13108] <= 1'b1;
startscreen[13125] <= 1'b1;
startscreen[13126] <= 1'b1;
startscreen[13127] <= 1'b1;
startscreen[13129] <= 1'b1;
startscreen[13165] <= 1'b1;
startscreen[13167] <= 1'b1;
startscreen[13174] <= 1'b1;
startscreen[13175] <= 1'b1;
startscreen[13176] <= 1'b1;
startscreen[13177] <= 1'b1;
startscreen[13192] <= 1'b1;
startscreen[13194] <= 1'b1;
startscreen[13195] <= 1'b1;
startscreen[13201] <= 1'b1;
startscreen[13203] <= 1'b1;
startscreen[13204] <= 1'b1;
startscreen[13216] <= 1'b1;
startscreen[13217] <= 1'b1;
startscreen[13218] <= 1'b1;
startscreen[13219] <= 1'b1;
startscreen[13225] <= 1'b1;
startscreen[13227] <= 1'b1;
startscreen[13228] <= 1'b1;
startscreen[13248] <= 1'b1;
startscreen[13250] <= 1'b1;
startscreen[13289] <= 1'b1;
startscreen[13291] <= 1'b1;
startscreen[13292] <= 1'b1;
startscreen[13302] <= 1'b1;
startscreen[13303] <= 1'b1;
startscreen[13304] <= 1'b1;
startscreen[13305] <= 1'b1;
startscreen[13322] <= 1'b1;
startscreen[13323] <= 1'b1;
startscreen[13324] <= 1'b1;
startscreen[13325] <= 1'b1;
startscreen[13360] <= 1'b1;
startscreen[13361] <= 1'b1;
startscreen[13362] <= 1'b1;
startscreen[13363] <= 1'b1;
startscreen[13370] <= 1'b1;
startscreen[13371] <= 1'b1;
startscreen[13372] <= 1'b1;
startscreen[13373] <= 1'b1;
startscreen[13383] <= 1'b1;
startscreen[13385] <= 1'b1;
startscreen[13386] <= 1'b1;
startscreen[13387] <= 1'b1;
startscreen[13398] <= 1'b1;
startscreen[13399] <= 1'b1;
startscreen[13400] <= 1'b1;
startscreen[13401] <= 1'b1;
startscreen[13402] <= 1'b1;
startscreen[13410] <= 1'b1;
startscreen[13412] <= 1'b1;
startscreen[13413] <= 1'b1;
startscreen[13427] <= 1'b1;
startscreen[13428] <= 1'b1;
startscreen[13430] <= 1'b1;
startscreen[13447] <= 1'b1;
startscreen[13448] <= 1'b1;
startscreen[13449] <= 1'b1;
startscreen[13450] <= 1'b1;
startscreen[13473] <= 1'b1;
startscreen[13474] <= 1'b1;
startscreen[13475] <= 1'b1;
startscreen[13476] <= 1'b1;
startscreen[13489] <= 1'b1;
startscreen[13490] <= 1'b1;
startscreen[13491] <= 1'b1;
startscreen[13492] <= 1'b1;
startscreen[13526] <= 1'b1;
startscreen[13527] <= 1'b1;
startscreen[13528] <= 1'b1;
startscreen[13529] <= 1'b1;
startscreen[13546] <= 1'b1;
startscreen[13547] <= 1'b1;
startscreen[13548] <= 1'b1;
startscreen[13549] <= 1'b1;
startscreen[13586] <= 1'b1;
startscreen[13587] <= 1'b1;
startscreen[13594] <= 1'b1;
startscreen[13595] <= 1'b1;
startscreen[13597] <= 1'b1;
startscreen[13613] <= 1'b1;
startscreen[13614] <= 1'b1;
startscreen[13615] <= 1'b1;
startscreen[13621] <= 1'b1;
startscreen[13622] <= 1'b1;
startscreen[13624] <= 1'b1;
startscreen[13636] <= 1'b1;
startscreen[13637] <= 1'b1;
startscreen[13639] <= 1'b1;
startscreen[13645] <= 1'b1;
startscreen[13646] <= 1'b1;
startscreen[13648] <= 1'b1;
startscreen[13649] <= 1'b1;
startscreen[13668] <= 1'b1;
startscreen[13669] <= 1'b1;
startscreen[13671] <= 1'b1;
startscreen[13709] <= 1'b1;
startscreen[13712] <= 1'b1;
startscreen[13723] <= 1'b1;
startscreen[13725] <= 1'b1;
startscreen[13726] <= 1'b1;
startscreen[13741] <= 1'b1;
startscreen[13742] <= 1'b1;
startscreen[13743] <= 1'b1;
startscreen[13744] <= 1'b1;
startscreen[13780] <= 1'b1;
startscreen[13781] <= 1'b1;
startscreen[13782] <= 1'b1;
startscreen[13783] <= 1'b1;
startscreen[13790] <= 1'b1;
startscreen[13792] <= 1'b1;
startscreen[13793] <= 1'b1;
startscreen[13803] <= 1'b1;
startscreen[13804] <= 1'b1;
startscreen[13806] <= 1'b1;
startscreen[13818] <= 1'b1;
startscreen[13819] <= 1'b1;
startscreen[13820] <= 1'b1;
startscreen[13821] <= 1'b1;
startscreen[13822] <= 1'b1;
startscreen[13830] <= 1'b1;
startscreen[13832] <= 1'b1;
startscreen[13833] <= 1'b1;
startscreen[13847] <= 1'b1;
startscreen[13848] <= 1'b1;
startscreen[13850] <= 1'b1;
startscreen[13867] <= 1'b1;
startscreen[13868] <= 1'b1;
startscreen[13869] <= 1'b1;
startscreen[13870] <= 1'b1;
startscreen[13893] <= 1'b1;
startscreen[13894] <= 1'b1;
startscreen[13895] <= 1'b1;
startscreen[13896] <= 1'b1;
startscreen[13909] <= 1'b1;
startscreen[13912] <= 1'b1;
startscreen[13913] <= 1'b1;
startscreen[13946] <= 1'b1;
startscreen[13948] <= 1'b1;
startscreen[13949] <= 1'b1;
startscreen[13966] <= 1'b1;
startscreen[13969] <= 1'b1;
startscreen[13987] <= 1'b1;
startscreen[13988] <= 1'b1;
startscreen[14004] <= 1'b1;
startscreen[14005] <= 1'b1;
startscreen[14007] <= 1'b1;
startscreen[14014] <= 1'b1;
startscreen[14015] <= 1'b1;
startscreen[14016] <= 1'b1;
startscreen[14017] <= 1'b1;
startscreen[14018] <= 1'b1;
startscreen[14031] <= 1'b1;
startscreen[14032] <= 1'b1;
startscreen[14033] <= 1'b1;
startscreen[14034] <= 1'b1;
startscreen[14041] <= 1'b1;
startscreen[14044] <= 1'b1;
startscreen[14055] <= 1'b1;
startscreen[14056] <= 1'b1;
startscreen[14058] <= 1'b1;
startscreen[14059] <= 1'b1;
startscreen[14066] <= 1'b1;
startscreen[14067] <= 1'b1;
startscreen[14068] <= 1'b1;
startscreen[14069] <= 1'b1;
startscreen[14070] <= 1'b1;
startscreen[14088] <= 1'b1;
startscreen[14089] <= 1'b1;
startscreen[14092] <= 1'b1;
startscreen[14130] <= 1'b1;
startscreen[14131] <= 1'b1;
startscreen[14132] <= 1'b1;
startscreen[14143] <= 1'b1;
startscreen[14144] <= 1'b1;
startscreen[14145] <= 1'b1;
startscreen[14146] <= 1'b1;
startscreen[14160] <= 1'b1;
startscreen[14161] <= 1'b1;
startscreen[14163] <= 1'b1;
startscreen[14164] <= 1'b1;
startscreen[14183] <= 1'b1;
startscreen[14184] <= 1'b1;
startscreen[14200] <= 1'b1;
startscreen[14201] <= 1'b1;
startscreen[14202] <= 1'b1;
startscreen[14203] <= 1'b1;
startscreen[14210] <= 1'b1;
startscreen[14211] <= 1'b1;
startscreen[14213] <= 1'b1;
startscreen[14223] <= 1'b1;
startscreen[14224] <= 1'b1;
startscreen[14225] <= 1'b1;
startscreen[14226] <= 1'b1;
startscreen[14238] <= 1'b1;
startscreen[14239] <= 1'b1;
startscreen[14240] <= 1'b1;
startscreen[14241] <= 1'b1;
startscreen[14242] <= 1'b1;
startscreen[14250] <= 1'b1;
startscreen[14252] <= 1'b1;
startscreen[14253] <= 1'b1;
startscreen[14267] <= 1'b1;
startscreen[14268] <= 1'b1;
startscreen[14287] <= 1'b1;
startscreen[14288] <= 1'b1;
startscreen[14289] <= 1'b1;
startscreen[14290] <= 1'b1;
startscreen[14313] <= 1'b1;
startscreen[14314] <= 1'b1;
startscreen[14315] <= 1'b1;
startscreen[14316] <= 1'b1;
startscreen[14332] <= 1'b1;
startscreen[14333] <= 1'b1;
startscreen[14334] <= 1'b1;
startscreen[14346] <= 1'b1;
startscreen[14347] <= 1'b1;
startscreen[14367] <= 1'b1;
startscreen[14368] <= 1'b1;
startscreen[14369] <= 1'b1;
startscreen[14386] <= 1'b1;
startscreen[14387] <= 1'b1;
startscreen[14389] <= 1'b1;
startscreen[14407] <= 1'b1;
startscreen[14408] <= 1'b1;
startscreen[14409] <= 1'b1;
startscreen[14423] <= 1'b1;
startscreen[14424] <= 1'b1;
startscreen[14427] <= 1'b1;
startscreen[14434] <= 1'b1;
startscreen[14435] <= 1'b1;
startscreen[14436] <= 1'b1;
startscreen[14437] <= 1'b1;
startscreen[14438] <= 1'b1;
startscreen[14439] <= 1'b1;
startscreen[14450] <= 1'b1;
startscreen[14451] <= 1'b1;
startscreen[14452] <= 1'b1;
startscreen[14454] <= 1'b1;
startscreen[14461] <= 1'b1;
startscreen[14462] <= 1'b1;
startscreen[14464] <= 1'b1;
startscreen[14474] <= 1'b1;
startscreen[14475] <= 1'b1;
startscreen[14476] <= 1'b1;
startscreen[14478] <= 1'b1;
startscreen[14479] <= 1'b1;
startscreen[14487] <= 1'b1;
startscreen[14488] <= 1'b1;
startscreen[14489] <= 1'b1;
startscreen[14490] <= 1'b1;
startscreen[14491] <= 1'b1;
startscreen[14509] <= 1'b1;
startscreen[14510] <= 1'b1;
startscreen[14511] <= 1'b1;
startscreen[14512] <= 1'b1;
startscreen[14525] <= 1'b1;
startscreen[14526] <= 1'b1;
startscreen[14549] <= 1'b1;
startscreen[14552] <= 1'b1;
startscreen[14564] <= 1'b1;
startscreen[14565] <= 1'b1;
startscreen[14566] <= 1'b1;
startscreen[14567] <= 1'b1;
startscreen[14580] <= 1'b1;
startscreen[14581] <= 1'b1;
startscreen[14582] <= 1'b1;
startscreen[14583] <= 1'b1;
startscreen[14603] <= 1'b1;
startscreen[14604] <= 1'b1;
startscreen[14605] <= 1'b1;
startscreen[14619] <= 1'b1;
startscreen[14620] <= 1'b1;
startscreen[14621] <= 1'b1;
startscreen[14622] <= 1'b1;
startscreen[14623] <= 1'b1;
startscreen[14630] <= 1'b1;
startscreen[14631] <= 1'b1;
startscreen[14632] <= 1'b1;
startscreen[14633] <= 1'b1;
startscreen[14643] <= 1'b1;
startscreen[14644] <= 1'b1;
startscreen[14646] <= 1'b1;
startscreen[14647] <= 1'b1;
startscreen[14657] <= 1'b1;
startscreen[14658] <= 1'b1;
startscreen[14659] <= 1'b1;
startscreen[14660] <= 1'b1;
startscreen[14661] <= 1'b1;
startscreen[14662] <= 1'b1;
startscreen[14670] <= 1'b1;
startscreen[14672] <= 1'b1;
startscreen[14673] <= 1'b1;
startscreen[14687] <= 1'b1;
startscreen[14688] <= 1'b1;
startscreen[14689] <= 1'b1;
startscreen[14690] <= 1'b1;
startscreen[14707] <= 1'b1;
startscreen[14708] <= 1'b1;
startscreen[14709] <= 1'b1;
startscreen[14710] <= 1'b1;
startscreen[14733] <= 1'b1;
startscreen[14734] <= 1'b1;
startscreen[14735] <= 1'b1;
startscreen[14736] <= 1'b1;
startscreen[14750] <= 1'b1;
startscreen[14751] <= 1'b1;
startscreen[14752] <= 1'b1;
startscreen[14754] <= 1'b1;
startscreen[14755] <= 1'b1;
startscreen[14765] <= 1'b1;
startscreen[14767] <= 1'b1;
startscreen[14773] <= 1'b1;
startscreen[14774] <= 1'b1;
startscreen[14785] <= 1'b1;
startscreen[14786] <= 1'b1;
startscreen[14788] <= 1'b1;
startscreen[14794] <= 1'b1;
startscreen[14795] <= 1'b1;
startscreen[14805] <= 1'b1;
startscreen[14806] <= 1'b1;
startscreen[14807] <= 1'b1;
startscreen[14808] <= 1'b1;
startscreen[14827] <= 1'b1;
startscreen[14828] <= 1'b1;
startscreen[14829] <= 1'b1;
startscreen[14830] <= 1'b1;
startscreen[14831] <= 1'b1;
startscreen[14842] <= 1'b1;
startscreen[14843] <= 1'b1;
startscreen[14844] <= 1'b1;
startscreen[14846] <= 1'b1;
startscreen[14854] <= 1'b1;
startscreen[14855] <= 1'b1;
startscreen[14857] <= 1'b1;
startscreen[14859] <= 1'b1;
startscreen[14860] <= 1'b1;
startscreen[14869] <= 1'b1;
startscreen[14870] <= 1'b1;
startscreen[14872] <= 1'b1;
startscreen[14873] <= 1'b1;
startscreen[14881] <= 1'b1;
startscreen[14882] <= 1'b1;
startscreen[14883] <= 1'b1;
startscreen[14884] <= 1'b1;
startscreen[14885] <= 1'b1;
startscreen[14893] <= 1'b1;
startscreen[14894] <= 1'b1;
startscreen[14896] <= 1'b1;
startscreen[14897] <= 1'b1;
startscreen[14899] <= 1'b1;
startscreen[14907] <= 1'b1;
startscreen[14908] <= 1'b1;
startscreen[14909] <= 1'b1;
startscreen[14911] <= 1'b1;
startscreen[14912] <= 1'b1;
startscreen[14922] <= 1'b1;
startscreen[14923] <= 1'b1;
startscreen[14929] <= 1'b1;
startscreen[14930] <= 1'b1;
startscreen[14931] <= 1'b1;
startscreen[14932] <= 1'b1;
startscreen[14933] <= 1'b1;
startscreen[14934] <= 1'b1;
startscreen[14944] <= 1'b1;
startscreen[14945] <= 1'b1;
startscreen[14946] <= 1'b1;
startscreen[14969] <= 1'b1;
startscreen[14970] <= 1'b1;
startscreen[14972] <= 1'b1;
startscreen[14984] <= 1'b1;
startscreen[14985] <= 1'b1;
startscreen[14986] <= 1'b1;
startscreen[14987] <= 1'b1;
startscreen[14988] <= 1'b1;
startscreen[14999] <= 1'b1;
startscreen[15000] <= 1'b1;
startscreen[15001] <= 1'b1;
startscreen[15002] <= 1'b1;
startscreen[15023] <= 1'b1;
startscreen[15024] <= 1'b1;
startscreen[15025] <= 1'b1;
startscreen[15026] <= 1'b1;
startscreen[15027] <= 1'b1;
startscreen[15036] <= 1'b1;
startscreen[15037] <= 1'b1;
startscreen[15038] <= 1'b1;
startscreen[15039] <= 1'b1;
startscreen[15041] <= 1'b1;
startscreen[15042] <= 1'b1;
startscreen[15050] <= 1'b1;
startscreen[15051] <= 1'b1;
startscreen[15053] <= 1'b1;
startscreen[15054] <= 1'b1;
startscreen[15063] <= 1'b1;
startscreen[15064] <= 1'b1;
startscreen[15065] <= 1'b1;
startscreen[15066] <= 1'b1;
startscreen[15067] <= 1'b1;
startscreen[15068] <= 1'b1;
startscreen[15076] <= 1'b1;
startscreen[15077] <= 1'b1;
startscreen[15078] <= 1'b1;
startscreen[15080] <= 1'b1;
startscreen[15081] <= 1'b1;
startscreen[15082] <= 1'b1;
startscreen[15090] <= 1'b1;
startscreen[15092] <= 1'b1;
startscreen[15093] <= 1'b1;
startscreen[15108] <= 1'b1;
startscreen[15110] <= 1'b1;
startscreen[15111] <= 1'b1;
startscreen[15127] <= 1'b1;
startscreen[15128] <= 1'b1;
startscreen[15129] <= 1'b1;
startscreen[15130] <= 1'b1;
startscreen[15153] <= 1'b1;
startscreen[15154] <= 1'b1;
startscreen[15155] <= 1'b1;
startscreen[15156] <= 1'b1;
startscreen[15171] <= 1'b1;
startscreen[15172] <= 1'b1;
startscreen[15174] <= 1'b1;
startscreen[15175] <= 1'b1;
startscreen[15176] <= 1'b1;
startscreen[15177] <= 1'b1;
startscreen[15182] <= 1'b1;
startscreen[15183] <= 1'b1;
startscreen[15186] <= 1'b1;
startscreen[15187] <= 1'b1;
startscreen[15193] <= 1'b1;
startscreen[15194] <= 1'b1;
startscreen[15195] <= 1'b1;
startscreen[15196] <= 1'b1;
startscreen[15203] <= 1'b1;
startscreen[15205] <= 1'b1;
startscreen[15207] <= 1'b1;
startscreen[15214] <= 1'b1;
startscreen[15215] <= 1'b1;
startscreen[15216] <= 1'b1;
startscreen[15217] <= 1'b1;
startscreen[15223] <= 1'b1;
startscreen[15224] <= 1'b1;
startscreen[15226] <= 1'b1;
startscreen[15228] <= 1'b1;
startscreen[15247] <= 1'b1;
startscreen[15248] <= 1'b1;
startscreen[15249] <= 1'b1;
startscreen[15250] <= 1'b1;
startscreen[15252] <= 1'b1;
startscreen[15253] <= 1'b1;
startscreen[15254] <= 1'b1;
startscreen[15259] <= 1'b1;
startscreen[15260] <= 1'b1;
startscreen[15261] <= 1'b1;
startscreen[15264] <= 1'b1;
startscreen[15265] <= 1'b1;
startscreen[15274] <= 1'b1;
startscreen[15275] <= 1'b1;
startscreen[15276] <= 1'b1;
startscreen[15277] <= 1'b1;
startscreen[15279] <= 1'b1;
startscreen[15280] <= 1'b1;
startscreen[15281] <= 1'b1;
startscreen[15282] <= 1'b1;
startscreen[15287] <= 1'b1;
startscreen[15288] <= 1'b1;
startscreen[15289] <= 1'b1;
startscreen[15291] <= 1'b1;
startscreen[15292] <= 1'b1;
startscreen[15302] <= 1'b1;
startscreen[15303] <= 1'b1;
startscreen[15305] <= 1'b1;
startscreen[15306] <= 1'b1;
startscreen[15312] <= 1'b1;
startscreen[15313] <= 1'b1;
startscreen[15314] <= 1'b1;
startscreen[15315] <= 1'b1;
startscreen[15316] <= 1'b1;
startscreen[15318] <= 1'b1;
startscreen[15319] <= 1'b1;
startscreen[15328] <= 1'b1;
startscreen[15329] <= 1'b1;
startscreen[15331] <= 1'b1;
startscreen[15332] <= 1'b1;
startscreen[15333] <= 1'b1;
startscreen[15339] <= 1'b1;
startscreen[15340] <= 1'b1;
startscreen[15341] <= 1'b1;
startscreen[15342] <= 1'b1;
startscreen[15343] <= 1'b1;
startscreen[15350] <= 1'b1;
startscreen[15351] <= 1'b1;
startscreen[15352] <= 1'b1;
startscreen[15353] <= 1'b1;
startscreen[15354] <= 1'b1;
startscreen[15355] <= 1'b1;
startscreen[15356] <= 1'b1;
startscreen[15362] <= 1'b1;
startscreen[15363] <= 1'b1;
startscreen[15364] <= 1'b1;
startscreen[15365] <= 1'b1;
startscreen[15366] <= 1'b1;
startscreen[15389] <= 1'b1;
startscreen[15390] <= 1'b1;
startscreen[15392] <= 1'b1;
startscreen[15393] <= 1'b1;
startscreen[15394] <= 1'b1;
startscreen[15397] <= 1'b1;
startscreen[15398] <= 1'b1;
startscreen[15405] <= 1'b1;
startscreen[15406] <= 1'b1;
startscreen[15409] <= 1'b1;
startscreen[15410] <= 1'b1;
startscreen[15416] <= 1'b1;
startscreen[15417] <= 1'b1;
startscreen[15418] <= 1'b1;
startscreen[15419] <= 1'b1;
startscreen[15420] <= 1'b1;
startscreen[15421] <= 1'b1;
startscreen[15443] <= 1'b1;
startscreen[15444] <= 1'b1;
startscreen[15448] <= 1'b1;
startscreen[15449] <= 1'b1;
startscreen[15450] <= 1'b1;
startscreen[15451] <= 1'b1;
startscreen[15455] <= 1'b1;
startscreen[15456] <= 1'b1;
startscreen[15458] <= 1'b1;
startscreen[15461] <= 1'b1;
startscreen[15471] <= 1'b1;
startscreen[15473] <= 1'b1;
startscreen[15474] <= 1'b1;
startscreen[15475] <= 1'b1;
startscreen[15479] <= 1'b1;
startscreen[15480] <= 1'b1;
startscreen[15484] <= 1'b1;
startscreen[15485] <= 1'b1;
startscreen[15486] <= 1'b1;
startscreen[15487] <= 1'b1;
startscreen[15488] <= 1'b1;
startscreen[15489] <= 1'b1;
startscreen[15490] <= 1'b1;
startscreen[15493] <= 1'b1;
startscreen[15494] <= 1'b1;
startscreen[15495] <= 1'b1;
startscreen[15496] <= 1'b1;
startscreen[15497] <= 1'b1;
startscreen[15498] <= 1'b1;
startscreen[15499] <= 1'b1;
startscreen[15500] <= 1'b1;
startscreen[15501] <= 1'b1;
startscreen[15502] <= 1'b1;
startscreen[15510] <= 1'b1;
startscreen[15512] <= 1'b1;
startscreen[15513] <= 1'b1;
startscreen[15528] <= 1'b1;
startscreen[15529] <= 1'b1;
startscreen[15531] <= 1'b1;
startscreen[15532] <= 1'b1;
startscreen[15536] <= 1'b1;
startscreen[15537] <= 1'b1;
startscreen[15547] <= 1'b1;
startscreen[15548] <= 1'b1;
startscreen[15549] <= 1'b1;
startscreen[15550] <= 1'b1;
startscreen[15573] <= 1'b1;
startscreen[15574] <= 1'b1;
startscreen[15575] <= 1'b1;
startscreen[15576] <= 1'b1;
startscreen[15592] <= 1'b1;
startscreen[15593] <= 1'b1;
startscreen[15594] <= 1'b1;
startscreen[15596] <= 1'b1;
startscreen[15597] <= 1'b1;
startscreen[15599] <= 1'b1;
startscreen[15600] <= 1'b1;
startscreen[15602] <= 1'b1;
startscreen[15603] <= 1'b1;
startscreen[15605] <= 1'b1;
startscreen[15607] <= 1'b1;
startscreen[15613] <= 1'b1;
startscreen[15618] <= 1'b1;
startscreen[15619] <= 1'b1;
startscreen[15621] <= 1'b1;
startscreen[15625] <= 1'b1;
startscreen[15626] <= 1'b1;
startscreen[15634] <= 1'b1;
startscreen[15636] <= 1'b1;
startscreen[15639] <= 1'b1;
startscreen[15641] <= 1'b1;
startscreen[15643] <= 1'b1;
startscreen[15644] <= 1'b1;
startscreen[15646] <= 1'b1;
startscreen[15647] <= 1'b1;
startscreen[15667] <= 1'b1;
startscreen[15668] <= 1'b1;
startscreen[15669] <= 1'b1;
startscreen[15670] <= 1'b1;
startscreen[15672] <= 1'b1;
startscreen[15674] <= 1'b1;
startscreen[15677] <= 1'b1;
startscreen[15678] <= 1'b1;
startscreen[15679] <= 1'b1;
startscreen[15682] <= 1'b1;
startscreen[15683] <= 1'b1;
startscreen[15684] <= 1'b1;
startscreen[15694] <= 1'b1;
startscreen[15695] <= 1'b1;
startscreen[15697] <= 1'b1;
startscreen[15700] <= 1'b1;
startscreen[15701] <= 1'b1;
startscreen[15702] <= 1'b1;
startscreen[15704] <= 1'b1;
startscreen[15705] <= 1'b1;
startscreen[15707] <= 1'b1;
startscreen[15708] <= 1'b1;
startscreen[15709] <= 1'b1;
startscreen[15711] <= 1'b1;
startscreen[15722] <= 1'b1;
startscreen[15723] <= 1'b1;
startscreen[15724] <= 1'b1;
startscreen[15725] <= 1'b1;
startscreen[15727] <= 1'b1;
startscreen[15728] <= 1'b1;
startscreen[15729] <= 1'b1;
startscreen[15730] <= 1'b1;
startscreen[15731] <= 1'b1;
startscreen[15732] <= 1'b1;
startscreen[15733] <= 1'b1;
startscreen[15734] <= 1'b1;
startscreen[15736] <= 1'b1;
startscreen[15737] <= 1'b1;
startscreen[15739] <= 1'b1;
startscreen[15749] <= 1'b1;
startscreen[15750] <= 1'b1;
startscreen[15751] <= 1'b1;
startscreen[15752] <= 1'b1;
startscreen[15753] <= 1'b1;
startscreen[15754] <= 1'b1;
startscreen[15755] <= 1'b1;
startscreen[15756] <= 1'b1;
startscreen[15758] <= 1'b1;
startscreen[15759] <= 1'b1;
startscreen[15760] <= 1'b1;
startscreen[15762] <= 1'b1;
startscreen[15763] <= 1'b1;
startscreen[15771] <= 1'b1;
startscreen[15772] <= 1'b1;
startscreen[15773] <= 1'b1;
startscreen[15774] <= 1'b1;
startscreen[15776] <= 1'b1;
startscreen[15777] <= 1'b1;
startscreen[15778] <= 1'b1;
startscreen[15784] <= 1'b1;
startscreen[15785] <= 1'b1;
startscreen[15786] <= 1'b1;
startscreen[15810] <= 1'b1;
startscreen[15811] <= 1'b1;
startscreen[15812] <= 1'b1;
startscreen[15813] <= 1'b1;
startscreen[15814] <= 1'b1;
startscreen[15815] <= 1'b1;
startscreen[15816] <= 1'b1;
startscreen[15817] <= 1'b1;
startscreen[15818] <= 1'b1;
startscreen[15826] <= 1'b1;
startscreen[15827] <= 1'b1;
startscreen[15828] <= 1'b1;
startscreen[15830] <= 1'b1;
startscreen[15831] <= 1'b1;
startscreen[15832] <= 1'b1;
startscreen[15833] <= 1'b1;
startscreen[15836] <= 1'b1;
startscreen[15837] <= 1'b1;
startscreen[15838] <= 1'b1;
startscreen[15839] <= 1'b1;
startscreen[15840] <= 1'b1;
startscreen[15864] <= 1'b1;
startscreen[15865] <= 1'b1;
startscreen[15866] <= 1'b1;
startscreen[15867] <= 1'b1;
startscreen[15870] <= 1'b1;
startscreen[15871] <= 1'b1;
startscreen[15872] <= 1'b1;
startscreen[15873] <= 1'b1;
startscreen[15874] <= 1'b1;
startscreen[15875] <= 1'b1;
startscreen[15876] <= 1'b1;
startscreen[15877] <= 1'b1;
startscreen[15878] <= 1'b1;
startscreen[15879] <= 1'b1;
startscreen[15880] <= 1'b1;
startscreen[15881] <= 1'b1;
startscreen[15891] <= 1'b1;
startscreen[15892] <= 1'b1;
startscreen[15895] <= 1'b1;
startscreen[15896] <= 1'b1;
startscreen[15897] <= 1'b1;
startscreen[15898] <= 1'b1;
startscreen[15899] <= 1'b1;
startscreen[15900] <= 1'b1;
startscreen[15905] <= 1'b1;
startscreen[15906] <= 1'b1;
startscreen[15908] <= 1'b1;
startscreen[15909] <= 1'b1;
startscreen[15910] <= 1'b1;
startscreen[15911] <= 1'b1;
startscreen[15912] <= 1'b1;
startscreen[15913] <= 1'b1;
startscreen[15914] <= 1'b1;
startscreen[15915] <= 1'b1;
startscreen[15916] <= 1'b1;
startscreen[15917] <= 1'b1;
startscreen[15920] <= 1'b1;
startscreen[15921] <= 1'b1;
startscreen[15922] <= 1'b1;
startscreen[15930] <= 1'b1;
startscreen[15932] <= 1'b1;
startscreen[15933] <= 1'b1;
startscreen[15949] <= 1'b1;
startscreen[15950] <= 1'b1;
startscreen[15951] <= 1'b1;
startscreen[15952] <= 1'b1;
startscreen[15953] <= 1'b1;
startscreen[15954] <= 1'b1;
startscreen[15955] <= 1'b1;
startscreen[15956] <= 1'b1;
startscreen[15957] <= 1'b1;
startscreen[15967] <= 1'b1;
startscreen[15968] <= 1'b1;
startscreen[15969] <= 1'b1;
startscreen[15970] <= 1'b1;
startscreen[15993] <= 1'b1;
startscreen[15994] <= 1'b1;
startscreen[15995] <= 1'b1;
startscreen[15996] <= 1'b1;
startscreen[16013] <= 1'b1;
startscreen[16014] <= 1'b1;
startscreen[16015] <= 1'b1;
startscreen[16017] <= 1'b1;
startscreen[16018] <= 1'b1;
startscreen[16021] <= 1'b1;
startscreen[16022] <= 1'b1;
startscreen[16023] <= 1'b1;
startscreen[16024] <= 1'b1;
startscreen[16025] <= 1'b1;
startscreen[16033] <= 1'b1;
startscreen[16035] <= 1'b1;
startscreen[16037] <= 1'b1;
startscreen[16039] <= 1'b1;
startscreen[16040] <= 1'b1;
startscreen[16042] <= 1'b1;
startscreen[16043] <= 1'b1;
startscreen[16044] <= 1'b1;
startscreen[16045] <= 1'b1;
startscreen[16054] <= 1'b1;
startscreen[16056] <= 1'b1;
startscreen[16057] <= 1'b1;
startscreen[16058] <= 1'b1;
startscreen[16059] <= 1'b1;
startscreen[16060] <= 1'b1;
startscreen[16062] <= 1'b1;
startscreen[16063] <= 1'b1;
startscreen[16065] <= 1'b1;
startscreen[16066] <= 1'b1;
startscreen[16089] <= 1'b1;
startscreen[16090] <= 1'b1;
startscreen[16091] <= 1'b1;
startscreen[16092] <= 1'b1;
startscreen[16093] <= 1'b1;
startscreen[16094] <= 1'b1;
startscreen[16096] <= 1'b1;
startscreen[16097] <= 1'b1;
startscreen[16099] <= 1'b1;
startscreen[16100] <= 1'b1;
startscreen[16102] <= 1'b1;
startscreen[16103] <= 1'b1;
startscreen[16114] <= 1'b1;
startscreen[16116] <= 1'b1;
startscreen[16117] <= 1'b1;
startscreen[16121] <= 1'b1;
startscreen[16123] <= 1'b1;
startscreen[16124] <= 1'b1;
startscreen[16125] <= 1'b1;
startscreen[16126] <= 1'b1;
startscreen[16127] <= 1'b1;
startscreen[16128] <= 1'b1;
startscreen[16129] <= 1'b1;
startscreen[16130] <= 1'b1;
startscreen[16143] <= 1'b1;
startscreen[16144] <= 1'b1;
startscreen[16145] <= 1'b1;
startscreen[16146] <= 1'b1;
startscreen[16149] <= 1'b1;
startscreen[16150] <= 1'b1;
startscreen[16151] <= 1'b1;
startscreen[16152] <= 1'b1;
startscreen[16153] <= 1'b1;
startscreen[16156] <= 1'b1;
startscreen[16157] <= 1'b1;
startscreen[16159] <= 1'b1;
startscreen[16170] <= 1'b1;
startscreen[16171] <= 1'b1;
startscreen[16172] <= 1'b1;
startscreen[16174] <= 1'b1;
startscreen[16175] <= 1'b1;
startscreen[16176] <= 1'b1;
startscreen[16177] <= 1'b1;
startscreen[16178] <= 1'b1;
startscreen[16179] <= 1'b1;
startscreen[16180] <= 1'b1;
startscreen[16181] <= 1'b1;
startscreen[16182] <= 1'b1;
startscreen[16183] <= 1'b1;
startscreen[16192] <= 1'b1;
startscreen[16193] <= 1'b1;
startscreen[16194] <= 1'b1;
startscreen[16195] <= 1'b1;
startscreen[16197] <= 1'b1;
startscreen[16198] <= 1'b1;
startscreen[16199] <= 1'b1;
startscreen[16200] <= 1'b1;
startscreen[16201] <= 1'b1;
startscreen[16202] <= 1'b1;
startscreen[16203] <= 1'b1;
startscreen[16204] <= 1'b1;
startscreen[16205] <= 1'b1;
startscreen[16230] <= 1'b1;
startscreen[16231] <= 1'b1;
startscreen[16232] <= 1'b1;
startscreen[16234] <= 1'b1;
startscreen[16237] <= 1'b1;
startscreen[16238] <= 1'b1;
startscreen[16248] <= 1'b1;
startscreen[16249] <= 1'b1;
startscreen[16250] <= 1'b1;
startscreen[16251] <= 1'b1;
startscreen[16252] <= 1'b1;
startscreen[16253] <= 1'b1;
startscreen[16254] <= 1'b1;
startscreen[16255] <= 1'b1;
startscreen[16256] <= 1'b1;
startscreen[16257] <= 1'b1;
startscreen[16258] <= 1'b1;
startscreen[16259] <= 1'b1;
startscreen[16285] <= 1'b1;
startscreen[16286] <= 1'b1;
startscreen[16287] <= 1'b1;
startscreen[16288] <= 1'b1;
startscreen[16291] <= 1'b1;
startscreen[16294] <= 1'b1;
startscreen[16296] <= 1'b1;
startscreen[16297] <= 1'b1;
startscreen[16298] <= 1'b1;
startscreen[16299] <= 1'b1;
startscreen[16300] <= 1'b1;
startscreen[16312] <= 1'b1;
startscreen[16313] <= 1'b1;
startscreen[16314] <= 1'b1;
startscreen[16315] <= 1'b1;
startscreen[16316] <= 1'b1;
startscreen[16317] <= 1'b1;
startscreen[16318] <= 1'b1;
startscreen[16319] <= 1'b1;
startscreen[16320] <= 1'b1;
startscreen[16326] <= 1'b1;
startscreen[16327] <= 1'b1;
startscreen[16328] <= 1'b1;
startscreen[16331] <= 1'b1;
startscreen[16332] <= 1'b1;
startscreen[16333] <= 1'b1;
startscreen[16334] <= 1'b1;
startscreen[16335] <= 1'b1;
startscreen[16339] <= 1'b1;
startscreen[16340] <= 1'b1;
startscreen[16341] <= 1'b1;
startscreen[16342] <= 1'b1;
startscreen[16350] <= 1'b1;
startscreen[16352] <= 1'b1;
startscreen[16353] <= 1'b1;
startscreen[16369] <= 1'b1;
startscreen[16371] <= 1'b1;
startscreen[16372] <= 1'b1;
startscreen[16373] <= 1'b1;
startscreen[16374] <= 1'b1;
startscreen[16375] <= 1'b1;
startscreen[16376] <= 1'b1;
startscreen[16377] <= 1'b1;
startscreen[16387] <= 1'b1;
startscreen[16388] <= 1'b1;
startscreen[16389] <= 1'b1;
startscreen[16390] <= 1'b1;
startscreen[16413] <= 1'b1;
startscreen[16414] <= 1'b1;
startscreen[16415] <= 1'b1;
startscreen[16416] <= 1'b1;
startscreen[16435] <= 1'b1;
startscreen[16436] <= 1'b1;
startscreen[16437] <= 1'b1;
startscreen[16438] <= 1'b1;
startscreen[16439] <= 1'b1;
startscreen[16440] <= 1'b1;
startscreen[16441] <= 1'b1;
startscreen[16442] <= 1'b1;
startscreen[16443] <= 1'b1;
startscreen[16456] <= 1'b1;
startscreen[16457] <= 1'b1;
startscreen[16458] <= 1'b1;
startscreen[16459] <= 1'b1;
startscreen[16460] <= 1'b1;
startscreen[16461] <= 1'b1;
startscreen[16462] <= 1'b1;
startscreen[16477] <= 1'b1;
startscreen[16478] <= 1'b1;
startscreen[16479] <= 1'b1;
startscreen[16480] <= 1'b1;
startscreen[16481] <= 1'b1;
startscreen[16482] <= 1'b1;
startscreen[16483] <= 1'b1;
startscreen[16513] <= 1'b1;
startscreen[16514] <= 1'b1;
startscreen[16515] <= 1'b1;
startscreen[16516] <= 1'b1;
startscreen[16517] <= 1'b1;
startscreen[16518] <= 1'b1;
startscreen[16519] <= 1'b1;
startscreen[16520] <= 1'b1;
startscreen[16534] <= 1'b1;
startscreen[16535] <= 1'b1;
startscreen[16536] <= 1'b1;
startscreen[16537] <= 1'b1;
startscreen[16542] <= 1'b1;
startscreen[16543] <= 1'b1;
startscreen[16544] <= 1'b1;
startscreen[16545] <= 1'b1;
startscreen[16546] <= 1'b1;
startscreen[16547] <= 1'b1;
startscreen[16548] <= 1'b1;
startscreen[16565] <= 1'b1;
startscreen[16566] <= 1'b1;
startscreen[16567] <= 1'b1;
startscreen[16568] <= 1'b1;
startscreen[16569] <= 1'b1;
startscreen[16570] <= 1'b1;
startscreen[16571] <= 1'b1;
startscreen[16572] <= 1'b1;
startscreen[16576] <= 1'b1;
startscreen[16577] <= 1'b1;
startscreen[16578] <= 1'b1;
startscreen[16579] <= 1'b1;
startscreen[16592] <= 1'b1;
startscreen[16593] <= 1'b1;
startscreen[16594] <= 1'b1;
startscreen[16595] <= 1'b1;
startscreen[16596] <= 1'b1;
startscreen[16597] <= 1'b1;
startscreen[16598] <= 1'b1;
startscreen[16599] <= 1'b1;
startscreen[16600] <= 1'b1;
startscreen[16614] <= 1'b1;
startscreen[16615] <= 1'b1;
startscreen[16616] <= 1'b1;
startscreen[16617] <= 1'b1;
startscreen[16618] <= 1'b1;
startscreen[16619] <= 1'b1;
startscreen[16620] <= 1'b1;
startscreen[16621] <= 1'b1;
startscreen[16622] <= 1'b1;
startscreen[16623] <= 1'b1;
startscreen[16652] <= 1'b1;
startscreen[16653] <= 1'b1;
startscreen[16654] <= 1'b1;
startscreen[16655] <= 1'b1;
startscreen[16656] <= 1'b1;
startscreen[16657] <= 1'b1;
startscreen[16658] <= 1'b1;
startscreen[16670] <= 1'b1;
startscreen[16671] <= 1'b1;
startscreen[16672] <= 1'b1;
startscreen[16673] <= 1'b1;
startscreen[16674] <= 1'b1;
startscreen[16675] <= 1'b1;
startscreen[16676] <= 1'b1;
startscreen[16677] <= 1'b1;
startscreen[16708] <= 1'b1;
startscreen[16709] <= 1'b1;
startscreen[16710] <= 1'b1;
startscreen[16711] <= 1'b1;
startscreen[16712] <= 1'b1;
startscreen[16713] <= 1'b1;
startscreen[16714] <= 1'b1;
startscreen[16715] <= 1'b1;
startscreen[16716] <= 1'b1;
startscreen[16717] <= 1'b1;
startscreen[16733] <= 1'b1;
startscreen[16734] <= 1'b1;
startscreen[16735] <= 1'b1;
startscreen[16736] <= 1'b1;
startscreen[16737] <= 1'b1;
startscreen[16738] <= 1'b1;
startscreen[16739] <= 1'b1;
startscreen[16748] <= 1'b1;
startscreen[16749] <= 1'b1;
startscreen[16750] <= 1'b1;
startscreen[16751] <= 1'b1;
startscreen[16752] <= 1'b1;
startscreen[16753] <= 1'b1;
startscreen[16759] <= 1'b1;
startscreen[16760] <= 1'b1;
startscreen[16770] <= 1'b1;
startscreen[16772] <= 1'b1;
startscreen[16773] <= 1'b1;
startscreen[16791] <= 1'b1;
startscreen[16792] <= 1'b1;
startscreen[16793] <= 1'b1;
startscreen[16794] <= 1'b1;
startscreen[16795] <= 1'b1;
startscreen[16796] <= 1'b1;
startscreen[16954] <= 1'b1;
startscreen[16955] <= 1'b1;
startscreen[16956] <= 1'b1;
startscreen[16957] <= 1'b1;
startscreen[17374] <= 1'b1;
startscreen[17375] <= 1'b1;
startscreen[17376] <= 1'b1;
startscreen[17377] <= 1'b1;
startscreen[17794] <= 1'b1;
startscreen[17795] <= 1'b1;
startscreen[17796] <= 1'b1;
startscreen[17797] <= 1'b1;
startscreen[18214] <= 1'b1;
startscreen[18215] <= 1'b1;
startscreen[18216] <= 1'b1;
startscreen[18217] <= 1'b1;
startscreen[18634] <= 1'b1;
startscreen[18635] <= 1'b1;
startscreen[18637] <= 1'b1;
startscreen[19054] <= 1'b1;
startscreen[19055] <= 1'b1;
startscreen[19056] <= 1'b1;
startscreen[19057] <= 1'b1;
startscreen[19474] <= 1'b1;
startscreen[19475] <= 1'b1;
startscreen[19477] <= 1'b1;
startscreen[19894] <= 1'b1;
startscreen[19895] <= 1'b1;
startscreen[19896] <= 1'b1;
startscreen[19897] <= 1'b1;
startscreen[20314] <= 1'b1;
startscreen[20316] <= 1'b1;
startscreen[20317] <= 1'b1;
startscreen[20734] <= 1'b1;
startscreen[20735] <= 1'b1;
startscreen[20737] <= 1'b1;


	 end
	 else
		 startscreen <= 1'b0;
	 

	 end
endmodule