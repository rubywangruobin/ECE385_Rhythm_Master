module dropper_twenty_three(input Reset, frame_clk, 
						 input logic [7:0] keycode,keycode_second,
						 output [9:0] drop23X, drop23Y,
						 output [1599:0] arrow23,
						 output logic score23);
	logic [9:0] arrow_X_Pos, arrow_Y_Pos, arrow_Y_Motion;
	logic [11:0] counter;
    parameter [9:0] X_start=160;  // Center position on the X axis
    parameter [9:0] Y_start=100;  // Center position on the Y axis
    parameter [9:0] Y_Max=400;     // Bottommost point on the Y axis
	 logic finish_on;
	 enum logic [3:0] {Halted, Normal, End} State, Next_state;
	 
	 always_ff @ (posedge frame_clk )
    begin
		if(Reset)
		begin
			State <= Halted;
		end	
		else if(State == Halted)
		begin
			counter = 0;
			score23 = 0;
			arrow_Y_Motion = 0; 
			arrow_Y_Pos = Y_start;
			State <= Next_state;
		end
		else if(State == Normal)
			begin
				if(counter <1560)
					counter = counter + 1;
				else
					begin
						arrow_Y_Motion = 1;
						if ((arrow_Y_Pos + 40) >= Y_Max)
							score23 = 1'b0;	
						else if ((keycode == 8'h07|| keycode_second == 8'h07) & (arrow_Y_Pos + 40 >= 340) & (arrow_Y_Pos + 40 < 400))
							score23 = 1'b1;
						else
						begin
							arrow_Y_Pos = (arrow_Y_Pos + arrow_Y_Motion); 
							counter = counter + 1;
						end
					end
				State <= Next_state;
			end
		else
			State <= Next_state;
    end
	 
	 always_comb
	 begin
		Next_state = State;
		finish_on = 1'b0;
		arrow_X_Pos = X_start;
		unique case(State)
			Halted:
			begin
				finish_on = 1'b0;
				if(keycode == 8'h2c)
					Next_state = Normal;
			end
			Normal:
				begin
				if(counter < 1560)
				begin
					Next_state = Normal;
					end
				else
					begin
						if ( (arrow_Y_Pos + 40) >= Y_Max )  
							begin
									finish_on = 1'b1; 
									Next_state = End;
							end
						 else if ((keycode == 8'h07|| keycode_second == 8'h07) & (arrow_Y_Pos + 40 >= 340) & (arrow_Y_Pos + 40 < 400))
							begin
									finish_on = 1'b1;
									Next_state = End;
							end
						 else
							begin
								  Next_state = Normal;
							end
					end
				end
			End:
				begin
				finish_on = 1;
				if(keycode == 8'h01)
					Next_state = Halted;
				end
		endcase
					
	 end
    assign drop23X = arrow_X_Pos;
   
    assign drop23Y = arrow_Y_Pos;
	 always_comb
	 begin
	 arrow23 <= 1'b0;
	 if(finish_on == 0)
	 begin
	 arrow23[420] <= 1'b1;
arrow23[421] <= 1'b1;
arrow23[460] <= 1'b1;
arrow23[461] <= 1'b1;
arrow23[500] <= 1'b1;
arrow23[501] <= 1'b1;
arrow23[502] <= 1'b1;
arrow23[503] <= 1'b1;
arrow23[540] <= 1'b1;
arrow23[541] <= 1'b1;
arrow23[542] <= 1'b1;
arrow23[543] <= 1'b1;
arrow23[580] <= 1'b1;
arrow23[581] <= 1'b1;
arrow23[582] <= 1'b1;
arrow23[583] <= 1'b1;
arrow23[584] <= 1'b1;
arrow23[585] <= 1'b1;
arrow23[620] <= 1'b1;
arrow23[621] <= 1'b1;
arrow23[622] <= 1'b1;
arrow23[623] <= 1'b1;
arrow23[624] <= 1'b1;
arrow23[625] <= 1'b1;
arrow23[648] <= 1'b1;
arrow23[649] <= 1'b1;
arrow23[650] <= 1'b1;
arrow23[651] <= 1'b1;
arrow23[652] <= 1'b1;
arrow23[653] <= 1'b1;
arrow23[654] <= 1'b1;
arrow23[655] <= 1'b1;
arrow23[656] <= 1'b1;
arrow23[657] <= 1'b1;
arrow23[658] <= 1'b1;
arrow23[659] <= 1'b1;
arrow23[660] <= 1'b1;
arrow23[661] <= 1'b1;
arrow23[662] <= 1'b1;
arrow23[663] <= 1'b1;
arrow23[664] <= 1'b1;
arrow23[665] <= 1'b1;
arrow23[666] <= 1'b1;
arrow23[667] <= 1'b1;
arrow23[688] <= 1'b1;
arrow23[689] <= 1'b1;
arrow23[690] <= 1'b1;
arrow23[691] <= 1'b1;
arrow23[692] <= 1'b1;
arrow23[693] <= 1'b1;
arrow23[694] <= 1'b1;
arrow23[695] <= 1'b1;
arrow23[696] <= 1'b1;
arrow23[697] <= 1'b1;
arrow23[698] <= 1'b1;
arrow23[699] <= 1'b1;
arrow23[700] <= 1'b1;
arrow23[701] <= 1'b1;
arrow23[702] <= 1'b1;
arrow23[703] <= 1'b1;
arrow23[704] <= 1'b1;
arrow23[705] <= 1'b1;
arrow23[706] <= 1'b1;
arrow23[707] <= 1'b1;
arrow23[728] <= 1'b1;
arrow23[729] <= 1'b1;
arrow23[730] <= 1'b1;
arrow23[731] <= 1'b1;
arrow23[732] <= 1'b1;
arrow23[733] <= 1'b1;
arrow23[734] <= 1'b1;
arrow23[735] <= 1'b1;
arrow23[736] <= 1'b1;
arrow23[737] <= 1'b1;
arrow23[738] <= 1'b1;
arrow23[739] <= 1'b1;
arrow23[740] <= 1'b1;
arrow23[741] <= 1'b1;
arrow23[742] <= 1'b1;
arrow23[743] <= 1'b1;
arrow23[744] <= 1'b1;
arrow23[745] <= 1'b1;
arrow23[746] <= 1'b1;
arrow23[747] <= 1'b1;
arrow23[748] <= 1'b1;
arrow23[749] <= 1'b1;
arrow23[768] <= 1'b1;
arrow23[769] <= 1'b1;
arrow23[770] <= 1'b1;
arrow23[771] <= 1'b1;
arrow23[772] <= 1'b1;
arrow23[773] <= 1'b1;
arrow23[774] <= 1'b1;
arrow23[775] <= 1'b1;
arrow23[776] <= 1'b1;
arrow23[777] <= 1'b1;
arrow23[778] <= 1'b1;
arrow23[779] <= 1'b1;
arrow23[780] <= 1'b1;
arrow23[781] <= 1'b1;
arrow23[782] <= 1'b1;
arrow23[783] <= 1'b1;
arrow23[784] <= 1'b1;
arrow23[785] <= 1'b1;
arrow23[786] <= 1'b1;
arrow23[787] <= 1'b1;
arrow23[788] <= 1'b1;
arrow23[789] <= 1'b1;
arrow23[808] <= 1'b1;
arrow23[809] <= 1'b1;
arrow23[810] <= 1'b1;
arrow23[811] <= 1'b1;
arrow23[812] <= 1'b1;
arrow23[813] <= 1'b1;
arrow23[814] <= 1'b1;
arrow23[815] <= 1'b1;
arrow23[816] <= 1'b1;
arrow23[817] <= 1'b1;
arrow23[818] <= 1'b1;
arrow23[819] <= 1'b1;
arrow23[820] <= 1'b1;
arrow23[821] <= 1'b1;
arrow23[822] <= 1'b1;
arrow23[823] <= 1'b1;
arrow23[824] <= 1'b1;
arrow23[825] <= 1'b1;
arrow23[826] <= 1'b1;
arrow23[827] <= 1'b1;
arrow23[848] <= 1'b1;
arrow23[849] <= 1'b1;
arrow23[850] <= 1'b1;
arrow23[851] <= 1'b1;
arrow23[852] <= 1'b1;
arrow23[853] <= 1'b1;
arrow23[854] <= 1'b1;
arrow23[855] <= 1'b1;
arrow23[856] <= 1'b1;
arrow23[857] <= 1'b1;
arrow23[858] <= 1'b1;
arrow23[859] <= 1'b1;
arrow23[860] <= 1'b1;
arrow23[861] <= 1'b1;
arrow23[862] <= 1'b1;
arrow23[863] <= 1'b1;
arrow23[864] <= 1'b1;
arrow23[865] <= 1'b1;
arrow23[866] <= 1'b1;
arrow23[867] <= 1'b1;
arrow23[900] <= 1'b1;
arrow23[901] <= 1'b1;
arrow23[902] <= 1'b1;
arrow23[903] <= 1'b1;
arrow23[904] <= 1'b1;
arrow23[905] <= 1'b1;
arrow23[940] <= 1'b1;
arrow23[941] <= 1'b1;
arrow23[942] <= 1'b1;
arrow23[943] <= 1'b1;
arrow23[944] <= 1'b1;
arrow23[945] <= 1'b1;
arrow23[980] <= 1'b1;
arrow23[981] <= 1'b1;
arrow23[982] <= 1'b1;
arrow23[983] <= 1'b1;
arrow23[1020] <= 1'b1;
arrow23[1021] <= 1'b1;
arrow23[1022] <= 1'b1;
arrow23[1023] <= 1'b1;
arrow23[1060] <= 1'b1;
arrow23[1061] <= 1'b1;
arrow23[1100] <= 1'b1;
arrow23[1101] <= 1'b1;


	 end
   else
		 arrow23 <= 1'b0;
end
endmodule